magic
tech scmos
timestamp 1597918584
<< nwell >>
rect -30 61 60 95
<< ntransistor >>
rect -14 45 -12 48
rect 7 45 9 48
rect -28 7 -26 32
rect 3 29 5 32
rect 16 29 18 32
<< ptransistor >>
rect -14 70 -12 73
rect 7 70 9 73
rect 30 70 32 73
<< ndiffusion >>
rect -24 45 -22 48
rect -18 45 -14 48
rect -12 45 -4 48
rect 0 45 7 48
rect 9 45 13 48
rect 17 45 19 48
rect -37 11 -28 32
rect -37 7 -35 11
rect -31 7 -28 11
rect -26 28 -25 32
rect -5 29 -4 32
rect 0 29 3 32
rect 5 29 8 32
rect -26 7 -21 28
rect 12 29 16 32
rect 18 29 23 32
rect 27 29 28 32
<< pdiffusion >>
rect -24 70 -22 73
rect -18 70 -14 73
rect -12 70 -4 73
rect 0 70 7 73
rect 9 70 13 73
rect 17 70 19 73
rect 22 70 23 73
rect 27 70 30 73
rect 32 70 35 73
rect 39 70 40 73
<< ndcontact >>
rect -22 45 -18 49
rect -4 44 0 48
rect 13 45 17 49
rect -35 7 -31 11
rect -25 28 -21 32
rect -4 29 0 33
rect 8 28 12 32
rect 23 29 27 33
<< pdcontact >>
rect -22 69 -18 73
rect -4 70 0 74
rect 13 69 17 73
rect 23 69 27 73
rect 35 70 39 74
<< psubstratepcontact >>
rect -3 15 1 19
rect 5 15 9 19
rect 13 15 17 19
<< nsubstratencontact >>
rect -15 85 -11 89
rect -7 85 -3 89
rect 1 85 5 89
rect 9 85 13 89
rect 17 85 21 89
rect 25 85 29 89
rect 33 85 37 89
<< polysilicon >>
rect -14 73 -12 76
rect 7 73 9 76
rect 30 73 32 76
rect -14 65 -12 70
rect 7 65 9 70
rect 30 67 32 70
rect -14 48 -12 51
rect 7 48 9 51
rect -14 42 -12 45
rect 7 42 9 45
rect -28 32 -26 35
rect 3 32 5 35
rect 16 32 18 35
rect 3 26 5 29
rect 16 26 18 29
rect -28 4 -26 7
<< polycontact >>
rect 28 76 32 80
rect -14 61 -10 65
rect 5 61 9 65
rect -29 35 -25 39
rect 3 35 7 39
rect 14 35 18 39
rect 1 22 5 26
<< metal1 >>
rect -19 85 -15 89
rect -11 85 -7 89
rect -3 85 1 89
rect 5 85 9 89
rect 13 85 17 89
rect 21 85 25 89
rect 29 85 33 89
rect 37 85 43 89
rect -4 74 0 85
rect 13 76 28 80
rect 13 73 17 76
rect 35 74 39 85
rect -22 49 -18 69
rect -10 61 5 65
rect 13 49 17 69
rect -39 35 -29 39
rect -25 35 -13 39
rect -25 32 -21 35
rect -17 26 -13 35
rect -4 33 0 44
rect 7 35 14 39
rect 23 33 27 69
rect -17 22 1 26
rect 8 19 12 28
rect -35 3 -31 7
rect -7 3 -3 19
rect 1 15 5 19
rect 9 15 13 19
rect 17 15 22 19
rect -35 -1 -3 3
<< labels >>
rlabel metal1 -2 86 -2 86 1 Vdd!
rlabel metal1 -5 17 -5 17 1 gnd!
<< end >>
