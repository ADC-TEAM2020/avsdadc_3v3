magic
tech scmos
timestamp 1599430094
<< nwell >>
rect 222 106 229 108
rect 451 106 457 108
rect 679 106 685 108
rect 907 106 916 108
rect 216 100 233 106
rect 445 100 461 106
rect 673 100 689 106
rect 901 100 920 106
rect 222 71 229 100
rect 451 71 457 100
rect 679 71 685 100
rect 907 71 916 100
rect -2 -21 4 -19
rect 226 -21 232 -19
rect 454 -21 460 -19
rect 682 -21 688 -19
rect 910 -21 916 -19
rect -6 -27 10 -21
rect 222 -27 238 -21
rect 450 -27 466 -21
rect 678 -27 694 -21
rect 906 -27 922 -21
rect -2 -56 4 -27
rect 226 -56 232 -27
rect 454 -56 460 -27
rect 682 -53 688 -27
rect 910 -56 916 -27
rect -2 -147 4 -145
rect 226 -147 232 -145
rect 454 -147 460 -145
rect 682 -147 688 -145
rect -8 -153 8 -147
rect 220 -153 236 -147
rect 448 -153 464 -147
rect 676 -153 692 -147
rect -2 -182 4 -153
rect 226 -158 232 -153
rect 226 -174 234 -158
rect 226 -182 232 -174
rect 454 -182 460 -153
rect 682 -182 688 -153
rect 910 -182 916 -145
rect 919 -158 923 -155
rect 919 -166 923 -162
rect 919 -182 923 -171
rect -228 -302 -224 -265
rect -2 -302 4 -265
rect 226 -302 232 -265
rect 454 -302 460 -265
rect 682 -267 688 -265
rect 910 -267 916 -265
rect 678 -273 694 -267
rect 906 -273 922 -267
rect 678 -290 681 -282
rect 682 -290 688 -273
rect 678 -294 688 -290
rect 682 -302 688 -294
rect 905 -295 909 -291
rect 910 -302 916 -273
rect -236 -415 -232 -378
rect -231 -548 -183 -491
rect 237 -597 767 -527
rect -145 -701 -97 -651
rect 17 -679 96 -599
rect 102 -679 154 -599
<< ntransistor >>
rect 252 -521 254 -511
rect 272 -521 274 -515
rect 305 -521 307 -511
rect 325 -521 327 -515
rect 358 -521 360 -511
rect 378 -521 380 -515
rect 411 -521 413 -511
rect 431 -521 433 -515
rect 464 -521 466 -511
rect 484 -521 486 -515
rect 517 -521 519 -511
rect 537 -521 539 -515
rect 570 -521 572 -511
rect 590 -521 592 -515
rect 623 -521 625 -511
rect 643 -521 645 -515
rect 676 -521 678 -511
rect 696 -521 698 -515
rect 729 -521 731 -511
rect 749 -521 751 -515
rect -216 -590 -214 -570
rect -211 -590 -209 -570
rect -203 -590 -201 -580
rect -133 -642 -131 -632
rect -115 -642 -113 -632
rect 31 -712 33 -692
rect 52 -712 54 -692
rect 117 -707 119 -697
rect 138 -707 140 -697
rect 15 -785 17 -765
rect 47 -779 49 -759
rect 68 -779 70 -759
<< ptransistor >>
rect -216 -522 -214 -502
rect -208 -522 -206 -502
rect -200 -522 -198 -502
rect 252 -573 254 -533
rect 272 -573 274 -561
rect 305 -573 307 -533
rect 325 -573 327 -561
rect 358 -573 360 -533
rect 378 -573 380 -561
rect 411 -573 413 -533
rect 431 -573 433 -561
rect 464 -573 466 -533
rect 484 -573 486 -561
rect 517 -573 519 -533
rect 537 -573 539 -561
rect 570 -573 572 -533
rect 590 -573 592 -561
rect 623 -573 625 -533
rect 643 -573 645 -561
rect 676 -573 678 -533
rect 696 -573 698 -561
rect 729 -573 731 -533
rect 749 -573 751 -561
rect -133 -677 -131 -657
rect -115 -677 -113 -657
rect 31 -670 33 -650
rect 52 -670 54 -650
rect 80 -670 82 -610
rect 117 -672 119 -652
rect 138 -672 140 -652
<< ndiffusion >>
rect 251 -521 252 -511
rect 254 -521 255 -511
rect 271 -521 272 -515
rect 274 -521 275 -515
rect 304 -521 305 -511
rect 307 -521 308 -511
rect 324 -521 325 -515
rect 327 -521 328 -515
rect 357 -521 358 -511
rect 360 -521 361 -511
rect 377 -521 378 -515
rect 380 -521 381 -515
rect 410 -521 411 -511
rect 413 -521 414 -511
rect 430 -521 431 -515
rect 433 -521 434 -515
rect 463 -521 464 -511
rect 466 -521 467 -511
rect 483 -521 484 -515
rect 486 -521 487 -515
rect 516 -521 517 -511
rect 519 -521 520 -511
rect 536 -521 537 -515
rect 539 -521 540 -515
rect 569 -521 570 -511
rect 572 -521 573 -511
rect 589 -521 590 -515
rect 592 -521 593 -515
rect 622 -521 623 -511
rect 625 -521 626 -511
rect 642 -521 643 -515
rect 645 -521 646 -515
rect 675 -521 676 -511
rect 678 -521 679 -511
rect 695 -521 696 -515
rect 698 -521 699 -515
rect 728 -521 729 -511
rect 731 -521 732 -511
rect 748 -521 749 -515
rect 751 -521 752 -515
rect -217 -590 -216 -570
rect -214 -590 -211 -570
rect -209 -590 -208 -570
rect -204 -590 -203 -580
rect -201 -590 -200 -580
rect -134 -642 -133 -632
rect -131 -642 -130 -632
rect -116 -642 -115 -632
rect -113 -642 -112 -632
rect 23 -696 24 -692
rect 28 -696 31 -692
rect 23 -697 31 -696
rect 23 -701 24 -697
rect 28 -701 31 -697
rect 23 -702 31 -701
rect 23 -706 24 -702
rect 28 -706 31 -702
rect 23 -707 31 -706
rect 23 -711 24 -707
rect 28 -711 31 -707
rect 23 -712 31 -711
rect 33 -693 41 -692
rect 33 -697 36 -693
rect 40 -697 41 -693
rect 33 -698 41 -697
rect 33 -702 36 -698
rect 40 -702 41 -698
rect 33 -703 41 -702
rect 33 -707 36 -703
rect 40 -707 41 -703
rect 33 -708 41 -707
rect 33 -712 36 -708
rect 40 -712 41 -708
rect 44 -696 45 -692
rect 49 -696 52 -692
rect 44 -697 52 -696
rect 44 -701 45 -697
rect 49 -701 52 -697
rect 44 -702 52 -701
rect 44 -706 45 -702
rect 49 -706 52 -702
rect 44 -707 52 -706
rect 44 -711 45 -707
rect 49 -711 52 -707
rect 44 -712 52 -711
rect 54 -693 62 -692
rect 54 -697 57 -693
rect 61 -697 62 -693
rect 54 -698 62 -697
rect 54 -702 57 -698
rect 61 -702 62 -698
rect 54 -703 62 -702
rect 54 -707 57 -703
rect 61 -707 62 -703
rect 109 -701 110 -697
rect 114 -701 117 -697
rect 109 -702 117 -701
rect 109 -706 110 -702
rect 114 -706 117 -702
rect 109 -707 117 -706
rect 119 -698 127 -697
rect 119 -702 122 -698
rect 126 -702 127 -698
rect 119 -703 127 -702
rect 119 -707 122 -703
rect 126 -707 127 -703
rect 130 -701 131 -697
rect 135 -701 138 -697
rect 130 -702 138 -701
rect 130 -706 131 -702
rect 135 -706 138 -702
rect 130 -707 138 -706
rect 140 -698 148 -697
rect 140 -702 143 -698
rect 147 -702 148 -698
rect 140 -703 148 -702
rect 140 -707 143 -703
rect 147 -707 148 -703
rect 54 -708 62 -707
rect 54 -712 57 -708
rect 61 -712 62 -708
rect 39 -763 40 -759
rect 44 -763 47 -759
rect 39 -764 47 -763
rect 7 -769 8 -765
rect 12 -769 15 -765
rect 7 -770 15 -769
rect 7 -774 8 -770
rect 12 -774 15 -770
rect 7 -775 15 -774
rect 7 -779 8 -775
rect 12 -779 15 -775
rect 7 -780 15 -779
rect 7 -784 8 -780
rect 12 -784 15 -780
rect 7 -785 15 -784
rect 17 -766 25 -765
rect 17 -770 20 -766
rect 24 -770 25 -766
rect 17 -771 25 -770
rect 17 -775 20 -771
rect 24 -775 25 -771
rect 17 -776 25 -775
rect 17 -780 20 -776
rect 24 -780 25 -776
rect 39 -768 40 -764
rect 44 -768 47 -764
rect 39 -769 47 -768
rect 39 -773 40 -769
rect 44 -773 47 -769
rect 39 -774 47 -773
rect 39 -778 40 -774
rect 44 -778 47 -774
rect 39 -779 47 -778
rect 49 -760 57 -759
rect 49 -764 52 -760
rect 56 -764 57 -760
rect 49 -765 57 -764
rect 49 -769 52 -765
rect 56 -769 57 -765
rect 49 -770 57 -769
rect 49 -774 52 -770
rect 56 -774 57 -770
rect 49 -775 57 -774
rect 49 -779 52 -775
rect 56 -779 57 -775
rect 60 -763 61 -759
rect 65 -763 68 -759
rect 60 -764 68 -763
rect 60 -768 61 -764
rect 65 -768 68 -764
rect 60 -769 68 -768
rect 60 -773 61 -769
rect 65 -773 68 -769
rect 60 -774 68 -773
rect 60 -778 61 -774
rect 65 -778 68 -774
rect 60 -779 68 -778
rect 70 -760 78 -759
rect 70 -764 73 -760
rect 77 -764 78 -760
rect 70 -765 78 -764
rect 70 -769 73 -765
rect 77 -769 78 -765
rect 70 -770 78 -769
rect 70 -774 73 -770
rect 77 -774 78 -770
rect 70 -775 78 -774
rect 70 -779 73 -775
rect 77 -779 78 -775
rect 17 -781 25 -780
rect 17 -785 20 -781
rect 24 -785 25 -781
<< pdiffusion >>
rect -217 -522 -216 -502
rect -214 -522 -213 -502
rect -209 -522 -208 -502
rect -206 -522 -205 -502
rect -201 -522 -200 -502
rect -198 -522 -197 -502
rect 251 -539 252 -533
rect 246 -545 252 -539
rect 251 -551 252 -545
rect 246 -557 252 -551
rect 251 -563 252 -557
rect 246 -567 252 -563
rect 251 -573 252 -567
rect 254 -539 255 -533
rect 254 -545 260 -539
rect 254 -551 255 -545
rect 254 -557 260 -551
rect 254 -563 255 -557
rect 304 -539 305 -533
rect 299 -545 305 -539
rect 304 -551 305 -545
rect 299 -557 305 -551
rect 254 -567 260 -563
rect 254 -573 255 -567
rect 271 -566 272 -561
rect 266 -568 272 -566
rect 271 -573 272 -568
rect 274 -566 275 -561
rect 274 -568 280 -566
rect 274 -573 275 -568
rect 304 -563 305 -557
rect 299 -567 305 -563
rect 304 -573 305 -567
rect 307 -539 308 -533
rect 307 -545 313 -539
rect 307 -551 308 -545
rect 307 -557 313 -551
rect 307 -563 308 -557
rect 357 -539 358 -533
rect 352 -545 358 -539
rect 357 -551 358 -545
rect 352 -557 358 -551
rect 307 -567 313 -563
rect 307 -573 308 -567
rect 324 -566 325 -561
rect 319 -568 325 -566
rect 324 -573 325 -568
rect 327 -566 328 -561
rect 327 -568 333 -566
rect 327 -573 328 -568
rect 357 -563 358 -557
rect 352 -567 358 -563
rect 357 -573 358 -567
rect 360 -539 361 -533
rect 360 -545 366 -539
rect 360 -551 361 -545
rect 360 -557 366 -551
rect 360 -563 361 -557
rect 410 -539 411 -533
rect 405 -545 411 -539
rect 410 -551 411 -545
rect 405 -557 411 -551
rect 360 -567 366 -563
rect 360 -573 361 -567
rect 377 -566 378 -561
rect 372 -568 378 -566
rect 377 -573 378 -568
rect 380 -566 381 -561
rect 380 -568 386 -566
rect 380 -573 381 -568
rect 410 -563 411 -557
rect 405 -567 411 -563
rect 410 -573 411 -567
rect 413 -539 414 -533
rect 413 -545 419 -539
rect 413 -551 414 -545
rect 413 -557 419 -551
rect 413 -563 414 -557
rect 463 -539 464 -533
rect 458 -545 464 -539
rect 463 -551 464 -545
rect 458 -557 464 -551
rect 413 -567 419 -563
rect 413 -573 414 -567
rect 430 -566 431 -561
rect 425 -568 431 -566
rect 430 -573 431 -568
rect 433 -566 434 -561
rect 433 -568 439 -566
rect 433 -573 434 -568
rect 463 -563 464 -557
rect 458 -567 464 -563
rect 463 -573 464 -567
rect 466 -539 467 -533
rect 466 -545 472 -539
rect 466 -551 467 -545
rect 466 -557 472 -551
rect 466 -563 467 -557
rect 516 -539 517 -533
rect 511 -545 517 -539
rect 516 -551 517 -545
rect 511 -557 517 -551
rect 466 -567 472 -563
rect 466 -573 467 -567
rect 483 -566 484 -561
rect 478 -568 484 -566
rect 483 -573 484 -568
rect 486 -566 487 -561
rect 486 -568 492 -566
rect 486 -573 487 -568
rect 516 -563 517 -557
rect 511 -567 517 -563
rect 516 -573 517 -567
rect 519 -539 520 -533
rect 519 -545 525 -539
rect 519 -551 520 -545
rect 519 -557 525 -551
rect 519 -563 520 -557
rect 569 -539 570 -533
rect 564 -545 570 -539
rect 569 -551 570 -545
rect 564 -557 570 -551
rect 519 -567 525 -563
rect 519 -573 520 -567
rect 536 -566 537 -561
rect 531 -568 537 -566
rect 536 -573 537 -568
rect 539 -566 540 -561
rect 539 -568 545 -566
rect 539 -573 540 -568
rect 569 -563 570 -557
rect 564 -567 570 -563
rect 569 -573 570 -567
rect 572 -539 573 -533
rect 572 -545 578 -539
rect 572 -551 573 -545
rect 572 -557 578 -551
rect 572 -563 573 -557
rect 622 -539 623 -533
rect 617 -545 623 -539
rect 622 -551 623 -545
rect 617 -557 623 -551
rect 572 -567 578 -563
rect 572 -573 573 -567
rect 589 -566 590 -561
rect 584 -568 590 -566
rect 589 -573 590 -568
rect 592 -566 593 -561
rect 592 -568 598 -566
rect 592 -573 593 -568
rect 622 -563 623 -557
rect 617 -567 623 -563
rect 622 -573 623 -567
rect 625 -539 626 -533
rect 625 -545 631 -539
rect 625 -551 626 -545
rect 625 -557 631 -551
rect 625 -563 626 -557
rect 675 -539 676 -533
rect 670 -545 676 -539
rect 675 -551 676 -545
rect 670 -557 676 -551
rect 625 -567 631 -563
rect 625 -573 626 -567
rect 642 -566 643 -561
rect 637 -568 643 -566
rect 642 -573 643 -568
rect 645 -566 646 -561
rect 645 -568 651 -566
rect 645 -573 646 -568
rect 675 -563 676 -557
rect 670 -567 676 -563
rect 675 -573 676 -567
rect 678 -539 679 -533
rect 678 -545 684 -539
rect 678 -551 679 -545
rect 678 -557 684 -551
rect 678 -563 679 -557
rect 728 -539 729 -533
rect 723 -545 729 -539
rect 728 -551 729 -545
rect 723 -557 729 -551
rect 678 -567 684 -563
rect 678 -573 679 -567
rect 695 -566 696 -561
rect 690 -568 696 -566
rect 695 -573 696 -568
rect 698 -566 699 -561
rect 698 -568 704 -566
rect 698 -573 699 -568
rect 728 -563 729 -557
rect 723 -567 729 -563
rect 728 -573 729 -567
rect 731 -539 732 -533
rect 731 -545 737 -539
rect 731 -551 732 -545
rect 731 -557 737 -551
rect 731 -563 732 -557
rect 731 -567 737 -563
rect 731 -573 732 -567
rect 748 -566 749 -561
rect 743 -568 749 -566
rect 748 -573 749 -568
rect 751 -566 752 -561
rect 751 -568 757 -566
rect 751 -573 752 -568
rect -134 -662 -133 -657
rect -139 -665 -133 -662
rect -134 -670 -133 -665
rect -139 -672 -133 -670
rect -134 -677 -133 -672
rect -131 -662 -130 -657
rect -131 -665 -125 -662
rect -131 -670 -130 -665
rect -131 -672 -125 -670
rect -131 -677 -130 -672
rect -116 -662 -115 -657
rect -121 -665 -115 -662
rect -116 -670 -115 -665
rect -121 -672 -115 -670
rect -116 -677 -115 -672
rect -113 -662 -112 -657
rect -113 -665 -107 -662
rect -113 -670 -112 -665
rect -113 -672 -107 -670
rect -113 -677 -112 -672
rect 72 -611 80 -610
rect 72 -615 73 -611
rect 77 -615 80 -611
rect 72 -616 80 -615
rect 72 -620 73 -616
rect 77 -620 80 -616
rect 72 -621 80 -620
rect 72 -625 73 -621
rect 77 -625 80 -621
rect 72 -626 80 -625
rect 72 -630 73 -626
rect 77 -630 80 -626
rect 72 -631 80 -630
rect 72 -635 73 -631
rect 77 -635 80 -631
rect 72 -636 80 -635
rect 72 -640 73 -636
rect 77 -640 80 -636
rect 72 -641 80 -640
rect 72 -645 73 -641
rect 77 -645 80 -641
rect 72 -646 80 -645
rect 72 -650 73 -646
rect 77 -650 80 -646
rect 23 -651 31 -650
rect 23 -655 24 -651
rect 28 -655 31 -651
rect 23 -656 31 -655
rect 23 -660 24 -656
rect 28 -660 31 -656
rect 23 -661 31 -660
rect 23 -665 24 -661
rect 28 -665 31 -661
rect 23 -666 31 -665
rect 23 -670 24 -666
rect 28 -670 31 -666
rect 33 -654 36 -650
rect 40 -654 41 -650
rect 33 -655 41 -654
rect 33 -659 36 -655
rect 40 -659 41 -655
rect 33 -660 41 -659
rect 33 -664 36 -660
rect 40 -664 41 -660
rect 33 -665 41 -664
rect 33 -669 36 -665
rect 40 -669 41 -665
rect 33 -670 41 -669
rect 44 -651 52 -650
rect 44 -655 45 -651
rect 49 -655 52 -651
rect 44 -656 52 -655
rect 44 -660 45 -656
rect 49 -660 52 -656
rect 44 -661 52 -660
rect 44 -665 45 -661
rect 49 -665 52 -661
rect 44 -666 52 -665
rect 44 -670 45 -666
rect 49 -670 52 -666
rect 54 -654 57 -650
rect 61 -654 62 -650
rect 54 -655 62 -654
rect 54 -659 57 -655
rect 61 -659 62 -655
rect 54 -660 62 -659
rect 54 -664 57 -660
rect 61 -664 62 -660
rect 54 -665 62 -664
rect 54 -669 57 -665
rect 61 -669 62 -665
rect 54 -670 62 -669
rect 72 -651 80 -650
rect 72 -655 73 -651
rect 77 -655 80 -651
rect 72 -656 80 -655
rect 72 -660 73 -656
rect 77 -660 80 -656
rect 72 -661 80 -660
rect 72 -665 73 -661
rect 77 -665 80 -661
rect 72 -666 80 -665
rect 72 -670 73 -666
rect 77 -670 80 -666
rect 82 -614 85 -610
rect 89 -614 90 -610
rect 82 -615 90 -614
rect 82 -619 85 -615
rect 89 -619 90 -615
rect 82 -620 90 -619
rect 82 -624 85 -620
rect 89 -624 90 -620
rect 82 -625 90 -624
rect 82 -629 85 -625
rect 89 -629 90 -625
rect 82 -630 90 -629
rect 82 -634 85 -630
rect 89 -634 90 -630
rect 82 -635 90 -634
rect 82 -639 85 -635
rect 89 -639 90 -635
rect 82 -640 90 -639
rect 82 -644 85 -640
rect 89 -644 90 -640
rect 82 -645 90 -644
rect 82 -649 85 -645
rect 89 -649 90 -645
rect 82 -650 90 -649
rect 82 -654 85 -650
rect 89 -654 90 -650
rect 82 -655 90 -654
rect 82 -659 85 -655
rect 89 -659 90 -655
rect 82 -660 90 -659
rect 82 -664 85 -660
rect 89 -664 90 -660
rect 82 -665 90 -664
rect 82 -669 85 -665
rect 89 -669 90 -665
rect 82 -670 90 -669
rect 109 -653 117 -652
rect 109 -657 110 -653
rect 114 -657 117 -653
rect 109 -658 117 -657
rect 109 -662 110 -658
rect 114 -662 117 -658
rect 109 -663 117 -662
rect 109 -667 110 -663
rect 114 -667 117 -663
rect 109 -668 117 -667
rect 109 -672 110 -668
rect 114 -672 117 -668
rect 119 -656 122 -652
rect 126 -656 127 -652
rect 119 -657 127 -656
rect 119 -661 122 -657
rect 126 -661 127 -657
rect 119 -662 127 -661
rect 119 -666 122 -662
rect 126 -666 127 -662
rect 119 -667 127 -666
rect 119 -671 122 -667
rect 126 -671 127 -667
rect 119 -672 127 -671
rect 130 -653 138 -652
rect 130 -657 131 -653
rect 135 -657 138 -653
rect 130 -658 138 -657
rect 130 -662 131 -658
rect 135 -662 138 -658
rect 130 -663 138 -662
rect 130 -667 131 -663
rect 135 -667 138 -663
rect 130 -668 138 -667
rect 130 -672 131 -668
rect 135 -672 138 -668
rect 140 -656 143 -652
rect 147 -656 148 -652
rect 140 -657 148 -656
rect 140 -661 143 -657
rect 147 -661 148 -657
rect 140 -662 148 -661
rect 140 -666 143 -662
rect 147 -666 148 -662
rect 140 -667 148 -666
rect 140 -671 143 -667
rect 147 -671 148 -667
rect 140 -672 148 -671
<< ndcontact >>
rect 246 -521 251 -511
rect 255 -521 260 -511
rect 266 -521 271 -515
rect 275 -521 280 -515
rect 299 -521 304 -511
rect 308 -521 313 -511
rect 319 -521 324 -515
rect 328 -521 333 -515
rect 352 -521 357 -511
rect 361 -521 366 -511
rect 372 -521 377 -515
rect 381 -521 386 -515
rect 405 -521 410 -511
rect 414 -521 419 -511
rect 425 -521 430 -515
rect 434 -521 439 -515
rect 458 -521 463 -511
rect 467 -521 472 -511
rect 478 -521 483 -515
rect 487 -521 492 -515
rect 511 -521 516 -511
rect 520 -521 525 -511
rect 531 -521 536 -515
rect 540 -521 545 -515
rect 564 -521 569 -511
rect 573 -521 578 -511
rect 584 -521 589 -515
rect 593 -521 598 -515
rect 617 -521 622 -511
rect 626 -521 631 -511
rect 637 -521 642 -515
rect 646 -521 651 -515
rect 670 -521 675 -511
rect 679 -521 684 -511
rect 690 -521 695 -515
rect 699 -521 704 -515
rect 723 -521 728 -511
rect 732 -521 737 -511
rect 743 -521 748 -515
rect 752 -521 757 -515
rect -221 -590 -217 -570
rect -208 -590 -204 -570
rect -200 -590 -196 -580
rect -139 -642 -134 -632
rect -130 -642 -125 -632
rect -121 -642 -116 -632
rect -112 -642 -107 -632
rect 24 -696 28 -692
rect 24 -701 28 -697
rect 24 -706 28 -702
rect 24 -711 28 -707
rect 36 -697 40 -693
rect 36 -702 40 -698
rect 36 -707 40 -703
rect 36 -712 40 -708
rect 45 -696 49 -692
rect 45 -701 49 -697
rect 45 -706 49 -702
rect 45 -711 49 -707
rect 57 -697 61 -693
rect 57 -702 61 -698
rect 57 -707 61 -703
rect 110 -701 114 -697
rect 110 -706 114 -702
rect 122 -702 126 -698
rect 122 -707 126 -703
rect 131 -701 135 -697
rect 131 -706 135 -702
rect 143 -702 147 -698
rect 143 -707 147 -703
rect 57 -712 61 -708
rect 40 -763 44 -759
rect 8 -769 12 -765
rect 8 -774 12 -770
rect 8 -779 12 -775
rect 8 -784 12 -780
rect 20 -770 24 -766
rect 20 -775 24 -771
rect 20 -780 24 -776
rect 40 -768 44 -764
rect 40 -773 44 -769
rect 40 -778 44 -774
rect 52 -764 56 -760
rect 52 -769 56 -765
rect 52 -774 56 -770
rect 52 -779 56 -775
rect 61 -763 65 -759
rect 61 -768 65 -764
rect 61 -773 65 -769
rect 61 -778 65 -774
rect 73 -764 77 -760
rect 73 -769 77 -765
rect 73 -774 77 -770
rect 73 -779 77 -775
rect 20 -785 24 -781
<< pdcontact >>
rect -221 -522 -217 -502
rect -213 -522 -209 -502
rect -205 -522 -201 -502
rect -197 -522 -193 -502
rect 246 -539 251 -533
rect 246 -551 251 -545
rect 246 -563 251 -557
rect 246 -573 251 -567
rect 255 -539 260 -533
rect 255 -551 260 -545
rect 255 -563 260 -557
rect 299 -539 304 -533
rect 299 -551 304 -545
rect 255 -573 260 -567
rect 266 -566 271 -561
rect 266 -573 271 -568
rect 275 -566 280 -561
rect 275 -573 280 -568
rect 299 -563 304 -557
rect 299 -573 304 -567
rect 308 -539 313 -533
rect 308 -551 313 -545
rect 308 -563 313 -557
rect 352 -539 357 -533
rect 352 -551 357 -545
rect 308 -573 313 -567
rect 319 -566 324 -561
rect 319 -573 324 -568
rect 328 -566 333 -561
rect 328 -573 333 -568
rect 352 -563 357 -557
rect 352 -573 357 -567
rect 361 -539 366 -533
rect 361 -551 366 -545
rect 361 -563 366 -557
rect 405 -539 410 -533
rect 405 -551 410 -545
rect 361 -573 366 -567
rect 372 -566 377 -561
rect 372 -573 377 -568
rect 381 -566 386 -561
rect 381 -573 386 -568
rect 405 -563 410 -557
rect 405 -573 410 -567
rect 414 -539 419 -533
rect 414 -551 419 -545
rect 414 -563 419 -557
rect 458 -539 463 -533
rect 458 -551 463 -545
rect 414 -573 419 -567
rect 425 -566 430 -561
rect 425 -573 430 -568
rect 434 -566 439 -561
rect 434 -573 439 -568
rect 458 -563 463 -557
rect 458 -573 463 -567
rect 467 -539 472 -533
rect 467 -551 472 -545
rect 467 -563 472 -557
rect 511 -539 516 -533
rect 511 -551 516 -545
rect 467 -573 472 -567
rect 478 -566 483 -561
rect 478 -573 483 -568
rect 487 -566 492 -561
rect 487 -573 492 -568
rect 511 -563 516 -557
rect 511 -573 516 -567
rect 520 -539 525 -533
rect 520 -551 525 -545
rect 520 -563 525 -557
rect 564 -539 569 -533
rect 564 -551 569 -545
rect 520 -573 525 -567
rect 531 -566 536 -561
rect 531 -573 536 -568
rect 540 -566 545 -561
rect 540 -573 545 -568
rect 564 -563 569 -557
rect 564 -573 569 -567
rect 573 -539 578 -533
rect 573 -551 578 -545
rect 573 -563 578 -557
rect 617 -539 622 -533
rect 617 -551 622 -545
rect 573 -573 578 -567
rect 584 -566 589 -561
rect 584 -573 589 -568
rect 593 -566 598 -561
rect 593 -573 598 -568
rect 617 -563 622 -557
rect 617 -573 622 -567
rect 626 -539 631 -533
rect 626 -551 631 -545
rect 626 -563 631 -557
rect 670 -539 675 -533
rect 670 -551 675 -545
rect 626 -573 631 -567
rect 637 -566 642 -561
rect 637 -573 642 -568
rect 646 -566 651 -561
rect 646 -573 651 -568
rect 670 -563 675 -557
rect 670 -573 675 -567
rect 679 -539 684 -533
rect 679 -551 684 -545
rect 679 -563 684 -557
rect 723 -539 728 -533
rect 723 -551 728 -545
rect 679 -573 684 -567
rect 690 -566 695 -561
rect 690 -573 695 -568
rect 699 -566 704 -561
rect 699 -573 704 -568
rect 723 -563 728 -557
rect 723 -573 728 -567
rect 732 -539 737 -533
rect 732 -551 737 -545
rect 732 -563 737 -557
rect 732 -573 737 -567
rect 743 -566 748 -561
rect 743 -573 748 -568
rect 752 -566 757 -561
rect 752 -573 757 -568
rect -139 -662 -134 -657
rect -139 -670 -134 -665
rect -139 -677 -134 -672
rect -130 -662 -125 -657
rect -130 -670 -125 -665
rect -130 -677 -125 -672
rect -121 -662 -116 -657
rect -121 -670 -116 -665
rect -121 -677 -116 -672
rect -112 -662 -107 -657
rect -112 -670 -107 -665
rect -112 -677 -107 -672
rect 73 -615 77 -611
rect 73 -620 77 -616
rect 73 -625 77 -621
rect 73 -630 77 -626
rect 73 -635 77 -631
rect 73 -640 77 -636
rect 73 -645 77 -641
rect 73 -650 77 -646
rect 24 -655 28 -651
rect 24 -660 28 -656
rect 24 -665 28 -661
rect 24 -670 28 -666
rect 36 -654 40 -650
rect 36 -659 40 -655
rect 36 -664 40 -660
rect 36 -669 40 -665
rect 45 -655 49 -651
rect 45 -660 49 -656
rect 45 -665 49 -661
rect 45 -670 49 -666
rect 57 -654 61 -650
rect 57 -659 61 -655
rect 57 -664 61 -660
rect 57 -669 61 -665
rect 73 -655 77 -651
rect 73 -660 77 -656
rect 73 -665 77 -661
rect 73 -670 77 -666
rect 85 -614 89 -610
rect 85 -619 89 -615
rect 85 -624 89 -620
rect 85 -629 89 -625
rect 85 -634 89 -630
rect 85 -639 89 -635
rect 85 -644 89 -640
rect 85 -649 89 -645
rect 85 -654 89 -650
rect 85 -659 89 -655
rect 85 -664 89 -660
rect 85 -669 89 -665
rect 110 -657 114 -653
rect 110 -662 114 -658
rect 110 -667 114 -663
rect 110 -672 114 -668
rect 122 -656 126 -652
rect 122 -661 126 -657
rect 122 -666 126 -662
rect 122 -671 126 -667
rect 131 -657 135 -653
rect 131 -662 135 -658
rect 131 -667 135 -663
rect 131 -672 135 -668
rect 143 -656 147 -652
rect 143 -661 147 -657
rect 143 -666 147 -662
rect 143 -671 147 -667
<< psubstratepcontact >>
rect -254 -372 -250 -368
rect -241 -372 -237 -368
rect -228 -372 -224 -368
rect -236 -485 -232 -481
rect -222 -485 -218 -481
rect -207 -485 -203 -481
rect 240 -503 244 -497
rect 251 -503 255 -497
rect 263 -503 267 -497
rect 273 -503 277 -497
rect 282 -503 286 -497
rect 293 -503 297 -497
rect 304 -503 308 -497
rect 316 -503 320 -497
rect 326 -503 330 -497
rect 335 -503 339 -497
rect 346 -503 350 -497
rect 357 -503 361 -497
rect 369 -503 373 -497
rect 379 -503 383 -497
rect 388 -503 392 -497
rect 399 -503 403 -497
rect 410 -503 414 -497
rect 422 -503 426 -497
rect 432 -503 436 -497
rect 441 -503 445 -497
rect 452 -503 456 -497
rect 463 -503 467 -497
rect 475 -503 479 -497
rect 485 -503 489 -497
rect 494 -503 498 -497
rect 505 -503 509 -497
rect 516 -503 520 -497
rect 528 -503 532 -497
rect 538 -503 542 -497
rect 547 -503 551 -497
rect 558 -503 562 -497
rect 569 -503 573 -497
rect 581 -503 585 -497
rect 591 -503 595 -497
rect 600 -503 604 -497
rect 611 -503 615 -497
rect 622 -503 626 -497
rect 634 -503 638 -497
rect 644 -503 648 -497
rect 653 -503 657 -497
rect 664 -503 668 -497
rect 675 -503 679 -497
rect 687 -503 691 -497
rect 697 -503 701 -497
rect 706 -503 710 -497
rect 717 -503 721 -497
rect 728 -503 732 -497
rect 740 -503 744 -497
rect 750 -503 754 -497
rect 759 -503 763 -497
rect -225 -598 -221 -594
rect -209 -598 -205 -594
rect -140 -626 -136 -620
rect -132 -626 -128 -620
rect -124 -626 -120 -620
rect -116 -626 -112 -620
rect -108 -626 -104 -620
rect 1 -793 5 -789
rect 9 -793 13 -789
rect 17 -793 21 -789
rect 25 -793 29 -789
rect 33 -793 37 -789
rect 41 -793 45 -789
rect 49 -793 53 -789
rect 57 -793 61 -789
rect 65 -793 69 -789
rect 73 -793 77 -789
rect 81 -793 85 -789
rect 104 -793 108 -789
rect 112 -793 116 -789
rect 120 -793 124 -789
rect 129 -793 133 -789
rect 137 -793 141 -789
rect 145 -793 149 -789
<< nsubstratencontact >>
rect -257 -272 -253 -268
rect -244 -272 -240 -268
rect -229 -272 -225 -268
rect -29 -272 -25 -268
rect -15 -272 -11 -268
rect -2 -272 2 -268
rect 18 -272 22 -268
rect -237 -385 -233 -381
rect -222 -385 -218 -381
rect -206 -385 -202 -381
rect -225 -498 -221 -494
rect -209 -498 -205 -494
rect 240 -593 244 -587
rect 250 -593 254 -587
rect 259 -593 263 -587
rect 267 -593 271 -587
rect 275 -593 279 -587
rect 283 -593 287 -587
rect 293 -593 297 -587
rect 303 -593 307 -587
rect 312 -593 316 -587
rect 320 -593 324 -587
rect 328 -593 332 -587
rect 336 -593 340 -587
rect 346 -593 350 -587
rect 356 -593 360 -587
rect 365 -593 369 -587
rect 373 -593 377 -587
rect 381 -593 385 -587
rect 389 -593 393 -587
rect 399 -593 403 -587
rect 409 -593 413 -587
rect 418 -593 422 -587
rect 426 -593 430 -587
rect 434 -593 438 -587
rect 442 -593 446 -587
rect 452 -593 456 -587
rect 462 -593 466 -587
rect 471 -593 475 -587
rect 479 -593 483 -587
rect 487 -593 491 -587
rect 495 -593 499 -587
rect 505 -593 509 -587
rect 515 -593 519 -587
rect 524 -593 528 -587
rect 532 -593 536 -587
rect 540 -593 544 -587
rect 548 -593 552 -587
rect 558 -593 562 -587
rect 568 -593 572 -587
rect 577 -593 581 -587
rect 585 -593 589 -587
rect 593 -593 597 -587
rect 601 -593 605 -587
rect 611 -593 615 -587
rect 621 -593 625 -587
rect 630 -593 634 -587
rect 638 -593 642 -587
rect 646 -593 650 -587
rect 654 -593 658 -587
rect 664 -593 668 -587
rect 674 -593 678 -587
rect 683 -593 687 -587
rect 691 -593 695 -587
rect 699 -593 703 -587
rect 707 -593 711 -587
rect 717 -593 721 -587
rect 727 -593 731 -587
rect 736 -593 740 -587
rect 744 -593 748 -587
rect 752 -593 756 -587
rect 760 -593 764 -587
rect 24 -606 28 -602
rect 32 -606 36 -602
rect 40 -606 44 -602
rect 48 -606 52 -602
rect 56 -606 60 -602
rect 64 -606 68 -602
rect 72 -606 76 -602
rect 80 -606 84 -602
rect 88 -606 92 -602
rect 105 -606 109 -602
rect 113 -606 117 -602
rect 121 -606 125 -602
rect 130 -606 134 -602
rect 138 -606 142 -602
rect -138 -697 -134 -691
rect -130 -697 -126 -691
rect -120 -697 -116 -691
rect -112 -697 -108 -691
rect -104 -697 -100 -691
rect -13 -617 -1 -611
rect -13 -753 -1 -747
rect 308 -632 320 -626
rect 308 -716 320 -710
rect 348 -633 360 -627
rect 348 -717 360 -711
rect 368 -633 380 -627
rect 368 -717 380 -711
rect 388 -633 400 -627
rect 388 -717 400 -711
rect 428 -633 440 -627
rect 428 -717 440 -711
rect 448 -633 460 -627
rect 448 -717 460 -711
rect 468 -633 480 -627
rect 468 -717 480 -711
rect 508 -633 520 -627
rect 508 -717 520 -711
rect 528 -633 540 -627
rect 528 -717 540 -711
rect 548 -633 560 -627
rect 548 -717 560 -711
rect 588 -633 600 -627
rect 588 -717 600 -711
rect 608 -633 620 -627
rect 608 -717 620 -711
rect 628 -633 640 -627
rect 628 -717 640 -711
rect 668 -633 680 -627
rect 668 -717 680 -711
rect 688 -633 700 -627
rect 688 -717 700 -711
rect 308 -733 320 -727
rect 308 -817 320 -811
rect 328 -733 340 -727
rect 328 -817 340 -811
rect 348 -733 360 -727
rect 348 -817 360 -811
rect 388 -733 400 -727
rect 388 -817 400 -811
rect 408 -733 420 -727
rect 408 -817 420 -811
rect 428 -733 440 -727
rect 428 -817 440 -811
rect 468 -733 480 -727
rect 468 -817 480 -811
rect 488 -733 500 -727
rect 488 -817 500 -811
rect 508 -733 520 -727
rect 508 -817 520 -811
rect 548 -733 560 -727
rect 548 -817 560 -811
rect 568 -733 580 -727
rect 568 -817 580 -811
rect 588 -733 600 -727
rect 588 -817 600 -811
rect 628 -733 640 -727
rect 628 -817 640 -811
rect 648 -733 660 -727
rect 648 -817 660 -811
rect 668 -733 680 -727
rect 668 -817 680 -811
<< polysilicon >>
rect -216 -502 -214 -500
rect -208 -502 -206 -500
rect -200 -502 -198 -500
rect 252 -511 254 -508
rect 268 -509 272 -489
rect 321 -508 325 -489
rect 374 -508 378 -489
rect 427 -508 431 -489
rect 480 -508 484 -489
rect 533 -508 537 -488
rect 586 -508 590 -488
rect 639 -508 643 -488
rect 692 -508 696 -489
rect 745 -508 749 -488
rect 268 -513 274 -509
rect 305 -511 307 -508
rect 272 -515 274 -513
rect 321 -513 327 -508
rect 358 -511 360 -508
rect 325 -515 327 -513
rect 374 -513 380 -508
rect 411 -511 413 -508
rect 378 -515 380 -513
rect 427 -513 433 -508
rect 464 -511 466 -508
rect 431 -515 433 -513
rect 480 -513 486 -508
rect 517 -511 519 -508
rect 484 -515 486 -513
rect 533 -513 539 -508
rect 570 -511 572 -508
rect 537 -515 539 -513
rect 586 -513 592 -508
rect 623 -511 625 -508
rect 590 -515 592 -513
rect 639 -513 645 -508
rect 676 -511 678 -508
rect 643 -515 645 -513
rect 692 -513 698 -508
rect 729 -511 731 -508
rect 696 -515 698 -513
rect 745 -513 751 -508
rect 749 -515 751 -513
rect -216 -555 -214 -522
rect -208 -543 -206 -522
rect -217 -559 -214 -555
rect -208 -557 -206 -547
rect -216 -570 -214 -559
rect -211 -559 -206 -557
rect -211 -570 -209 -559
rect -200 -563 -198 -522
rect 252 -533 254 -521
rect -199 -566 -198 -563
rect -203 -580 -201 -567
rect 272 -561 274 -521
rect 305 -533 307 -521
rect 325 -561 327 -521
rect 358 -533 360 -521
rect 378 -561 380 -521
rect 411 -533 413 -521
rect 431 -561 433 -521
rect 464 -533 466 -521
rect 484 -561 486 -521
rect 517 -533 519 -521
rect 537 -561 539 -521
rect 570 -533 572 -521
rect 590 -561 592 -521
rect 623 -533 625 -521
rect 643 -561 645 -521
rect 676 -533 678 -521
rect 696 -561 698 -521
rect 729 -533 731 -521
rect 749 -561 751 -521
rect 252 -579 254 -573
rect 272 -576 274 -573
rect 305 -579 307 -573
rect 325 -576 327 -573
rect 358 -579 360 -573
rect 378 -576 380 -573
rect 411 -579 413 -573
rect 431 -576 433 -573
rect 464 -579 466 -573
rect 484 -576 486 -573
rect 517 -579 519 -573
rect 537 -576 539 -573
rect 570 -579 572 -573
rect 590 -576 592 -573
rect 623 -579 625 -573
rect 643 -576 645 -573
rect 676 -579 678 -573
rect 696 -576 698 -573
rect 729 -579 731 -573
rect 749 -576 751 -573
rect 252 -583 276 -579
rect 305 -583 329 -579
rect 358 -583 382 -579
rect 411 -583 435 -579
rect 464 -583 488 -579
rect 517 -583 541 -579
rect 570 -583 594 -579
rect 623 -583 647 -579
rect 676 -583 700 -579
rect 729 -583 753 -579
rect -216 -592 -214 -590
rect -211 -592 -209 -590
rect -203 -592 -201 -590
rect 80 -610 82 -607
rect -133 -630 -113 -628
rect -133 -632 -131 -630
rect -115 -632 -113 -630
rect -133 -651 -131 -642
rect -115 -645 -113 -642
rect -143 -656 -131 -651
rect -133 -657 -131 -656
rect -115 -657 -113 -655
rect -133 -680 -131 -677
rect -115 -683 -113 -677
rect -125 -687 -113 -683
rect 31 -650 33 -647
rect 52 -650 54 -647
rect 117 -652 119 -649
rect 138 -652 140 -649
rect 31 -675 33 -670
rect 52 -675 54 -670
rect 80 -678 82 -670
rect 31 -692 33 -689
rect 52 -692 54 -687
rect 117 -697 119 -672
rect 138 -697 140 -672
rect 117 -710 119 -707
rect 138 -710 140 -707
rect 31 -717 33 -712
rect 52 -715 54 -712
rect 47 -759 49 -748
rect 68 -759 70 -748
rect 15 -765 17 -762
rect 47 -782 49 -779
rect 68 -782 70 -779
rect 15 -788 17 -785
<< polycontact >>
rect 268 -489 272 -484
rect 321 -489 325 -484
rect 374 -489 378 -484
rect 427 -489 431 -484
rect 480 -489 484 -484
rect 533 -488 537 -483
rect 586 -488 590 -484
rect 639 -488 643 -484
rect 692 -489 696 -484
rect 745 -488 749 -483
rect -210 -547 -206 -543
rect -221 -559 -217 -555
rect -203 -567 -199 -563
rect 276 -583 280 -579
rect 329 -583 333 -579
rect 382 -583 386 -579
rect 435 -583 439 -579
rect 488 -583 492 -579
rect 541 -583 545 -579
rect 594 -583 598 -579
rect 647 -583 651 -579
rect 700 -583 704 -579
rect 753 -583 757 -579
rect -148 -656 -143 -651
rect -130 -687 -125 -683
rect 31 -679 35 -675
rect 50 -679 54 -675
rect 82 -678 86 -674
rect 50 -687 54 -683
rect 113 -693 117 -689
rect 134 -693 138 -689
rect 31 -721 35 -717
rect 47 -748 51 -744
rect 66 -748 70 -744
rect 15 -762 19 -758
<< metal1 >>
rect 216 100 233 106
rect 445 100 461 106
rect 673 100 689 106
rect 901 100 920 106
rect 1132 100 1157 106
rect 2 63 3 67
rect 445 63 460 67
rect 673 63 688 67
rect 902 63 919 67
rect 217 54 225 58
rect 446 54 453 58
rect 674 54 681 58
rect 902 54 909 58
rect 1133 54 1168 58
rect -19 50 3 54
rect -19 6 -15 50
rect 221 44 225 54
rect 449 44 453 54
rect 677 44 681 54
rect 905 44 909 54
rect 916 50 919 54
rect -10 40 3 44
rect 221 40 232 44
rect 453 40 460 44
rect 681 40 688 44
rect 909 40 919 44
rect -10 6 -6 40
rect 210 6 214 26
rect 441 6 445 9
rect 669 6 674 9
rect 897 7 898 11
rect 897 6 902 7
rect -19 0 3 6
rect 216 0 232 6
rect 445 0 460 6
rect 673 0 688 6
rect 901 0 919 6
rect -6 -27 10 -21
rect 222 -27 238 -21
rect 450 -27 466 -21
rect 678 -27 694 -21
rect 906 -27 922 -21
rect 1134 -27 1157 -21
rect -231 -73 -219 -69
rect 2 -73 9 -69
rect 230 -73 237 -69
rect 458 -73 465 -69
rect 686 -73 693 -69
rect -230 -186 -226 -73
rect 2 -83 6 -73
rect 230 -83 234 -73
rect 458 -83 462 -73
rect 686 -83 690 -73
rect 914 -83 918 -69
rect 1164 -83 1168 54
rect -5 -87 2 -83
rect 223 -87 234 -83
rect 451 -87 462 -83
rect 679 -87 690 -83
rect 907 -87 918 -83
rect 1135 -87 1164 -83
rect 230 -94 234 -87
rect 458 -95 462 -87
rect -13 -121 -9 -102
rect 215 -121 219 -102
rect 686 -95 690 -87
rect 905 -94 914 -90
rect 443 -121 447 -102
rect 671 -121 675 -103
rect 899 -121 903 -103
rect 1127 -108 1131 -103
rect 1130 -121 1131 -108
rect -5 -127 10 -121
rect 223 -127 238 -121
rect 451 -127 466 -121
rect 679 -127 694 -121
rect 907 -127 922 -121
rect 1135 -127 1149 -121
rect -8 -153 8 -147
rect 220 -153 236 -147
rect 448 -153 464 -147
rect 676 -153 692 -147
rect 904 -153 920 -147
rect 1132 -153 1157 -147
rect 918 -186 922 -183
rect -230 -190 -221 -186
rect 6 -190 7 -186
rect 234 -190 237 -186
rect 462 -190 463 -186
rect 690 -190 691 -186
rect 918 -190 919 -186
rect -7 -199 0 -195
rect 221 -199 228 -195
rect 449 -199 456 -195
rect 677 -199 684 -195
rect 905 -199 912 -195
rect 1132 -199 1152 -195
rect -220 -253 -216 -199
rect -4 -216 0 -199
rect 8 -203 10 -199
rect -4 -220 7 -216
rect 224 -220 228 -199
rect 232 -220 235 -216
rect 452 -220 456 -199
rect 460 -220 463 -216
rect 680 -220 684 -199
rect 694 -213 696 -209
rect 688 -220 691 -216
rect 908 -220 912 -199
rect 916 -220 919 -216
rect -8 -253 7 -247
rect 219 -253 235 -247
rect 447 -253 463 -247
rect 676 -253 691 -247
rect 903 -253 919 -247
rect -466 -273 -446 -267
rect -234 -268 -220 -267
rect -8 -268 10 -267
rect -234 -272 -229 -268
rect -225 -272 -220 -268
rect -8 -272 -2 -268
rect 2 -272 10 -268
rect -234 -273 -220 -272
rect -8 -273 10 -272
rect 222 -273 238 -267
rect 450 -273 466 -267
rect 678 -273 694 -267
rect 906 -273 922 -267
rect -466 -380 -461 -273
rect -447 -319 -444 -306
rect -221 -319 -218 -306
rect 221 -310 225 -302
rect 449 -310 453 -303
rect 677 -310 681 -303
rect 905 -310 909 -303
rect 1138 -310 1145 -306
rect -456 -323 -444 -319
rect -230 -323 -218 -319
rect 1 -319 9 -315
rect 230 -319 237 -315
rect 458 -319 465 -315
rect 686 -319 693 -315
rect 914 -319 920 -315
rect -456 -367 -452 -323
rect -230 -367 -226 -323
rect 1 -346 5 -319
rect 230 -336 234 -319
rect 458 -336 462 -319
rect 686 -336 690 -319
rect 914 -336 918 -319
rect 1135 -333 1140 -329
rect 1148 -336 1152 -199
rect 223 -340 237 -336
rect 451 -340 462 -336
rect 679 -340 690 -336
rect 907 -340 918 -336
rect 1135 -340 1167 -336
rect 1133 -367 1137 -361
rect -456 -373 -447 -367
rect -235 -368 -221 -367
rect -235 -372 -228 -368
rect -224 -372 -221 -368
rect -235 -373 -221 -372
rect -8 -373 13 -367
rect 223 -373 238 -367
rect 451 -373 466 -367
rect 679 -373 694 -367
rect 907 -373 922 -367
rect 1135 -373 1155 -367
rect -466 -386 -452 -380
rect -240 -381 -226 -380
rect -240 -385 -237 -381
rect -233 -385 -226 -381
rect -240 -386 -226 -385
rect -466 -493 -461 -386
rect -239 -423 -230 -419
rect -234 -480 -230 -423
rect -16 -432 -13 -419
rect -8 -432 -4 -373
rect 1163 -389 1167 -340
rect 1 -397 5 -391
rect 569 -393 959 -389
rect 1 -401 1167 -397
rect -16 -436 -4 -432
rect -8 -480 -4 -436
rect -239 -481 -226 -480
rect -239 -485 -236 -481
rect -232 -485 -226 -481
rect -239 -486 -226 -485
rect -13 -486 -4 -480
rect 219 -484 223 -401
rect 1159 -408 1167 -404
rect 321 -484 325 -465
rect -466 -499 -448 -493
rect -237 -494 -189 -493
rect -237 -498 -225 -494
rect -221 -498 -209 -494
rect -205 -498 -189 -494
rect -237 -499 -189 -498
rect -221 -502 -217 -499
rect -205 -502 -201 -499
rect -212 -525 -209 -522
rect -212 -528 -200 -525
rect -459 -536 -450 -532
rect -459 -593 -455 -536
rect -236 -545 -210 -541
rect -226 -559 -221 -555
rect -203 -563 -200 -528
rect -214 -566 -203 -563
rect -221 -570 -211 -566
rect -196 -566 -193 -522
rect -196 -577 -193 -570
rect -200 -580 -193 -577
rect -208 -593 -204 -590
rect -185 -593 -181 -486
rect 219 -489 268 -484
rect 374 -484 378 -465
rect 427 -484 431 -466
rect 480 -484 484 -414
rect 1159 -415 1167 -411
rect 1159 -422 1167 -418
rect 1159 -429 1167 -425
rect 1159 -436 1167 -432
rect 1159 -443 1167 -439
rect 1159 -450 1167 -446
rect 533 -483 537 -467
rect 586 -484 590 -455
rect 1159 -457 1167 -453
rect 1159 -464 1167 -460
rect 639 -484 643 -474
rect 692 -484 696 -471
rect 745 -483 749 -478
rect 237 -497 772 -496
rect 237 -503 240 -497
rect 244 -503 251 -497
rect 255 -503 263 -497
rect 267 -503 273 -497
rect 277 -503 282 -497
rect 286 -503 293 -497
rect 297 -503 304 -497
rect 308 -503 316 -497
rect 320 -503 326 -497
rect 330 -503 335 -497
rect 339 -503 346 -497
rect 350 -503 357 -497
rect 361 -503 369 -497
rect 373 -503 379 -497
rect 383 -503 388 -497
rect 392 -503 399 -497
rect 403 -503 410 -497
rect 414 -503 422 -497
rect 426 -503 432 -497
rect 436 -503 441 -497
rect 445 -503 452 -497
rect 456 -503 463 -497
rect 467 -503 475 -497
rect 479 -503 485 -497
rect 489 -503 494 -497
rect 498 -503 505 -497
rect 509 -503 516 -497
rect 520 -503 528 -497
rect 532 -503 538 -497
rect 542 -503 547 -497
rect 551 -503 558 -497
rect 562 -503 569 -497
rect 573 -503 581 -497
rect 585 -503 591 -497
rect 595 -503 600 -497
rect 604 -503 611 -497
rect 615 -503 622 -497
rect 626 -503 634 -497
rect 638 -503 644 -497
rect 648 -503 653 -497
rect 657 -503 664 -497
rect 668 -503 675 -497
rect 679 -503 687 -497
rect 691 -503 697 -497
rect 701 -503 706 -497
rect 710 -503 717 -497
rect 721 -503 728 -497
rect 732 -503 740 -497
rect 744 -503 750 -497
rect 754 -503 759 -497
rect 763 -503 772 -497
rect 237 -504 772 -503
rect 246 -511 251 -504
rect 266 -515 271 -504
rect 299 -511 304 -504
rect 319 -515 324 -504
rect 352 -511 357 -504
rect 372 -515 377 -504
rect 405 -511 410 -504
rect 425 -515 430 -504
rect 458 -511 463 -504
rect 478 -515 483 -504
rect 511 -511 516 -504
rect 531 -515 536 -504
rect 564 -511 569 -504
rect 584 -515 589 -504
rect 617 -511 622 -504
rect 637 -515 642 -504
rect 670 -511 675 -504
rect 690 -515 695 -504
rect 723 -511 728 -504
rect 743 -515 748 -504
rect 225 -533 231 -527
rect 246 -545 251 -539
rect 246 -557 251 -551
rect 246 -567 251 -563
rect 255 -533 260 -521
rect 255 -545 260 -539
rect 255 -557 260 -551
rect 275 -561 280 -521
rect 255 -567 260 -563
rect 266 -568 271 -566
rect 275 -568 280 -566
rect 299 -545 304 -539
rect 299 -557 304 -551
rect 299 -567 304 -563
rect 308 -533 313 -521
rect 308 -545 313 -539
rect 308 -557 313 -551
rect 328 -561 333 -521
rect 308 -567 313 -563
rect 319 -568 324 -566
rect 328 -568 333 -566
rect 352 -545 357 -539
rect 352 -557 357 -551
rect 352 -567 357 -563
rect 361 -533 366 -521
rect 361 -545 366 -539
rect 361 -557 366 -551
rect 381 -561 386 -521
rect 361 -567 366 -563
rect 372 -568 377 -566
rect 381 -568 386 -566
rect 405 -545 410 -539
rect 405 -557 410 -551
rect 405 -567 410 -563
rect 414 -533 419 -521
rect 414 -545 419 -539
rect 414 -557 419 -551
rect 434 -561 439 -521
rect 414 -567 419 -563
rect 425 -568 430 -566
rect 434 -568 439 -566
rect 458 -545 463 -539
rect 458 -557 463 -551
rect 458 -567 463 -563
rect 467 -533 472 -521
rect 467 -545 472 -539
rect 467 -557 472 -551
rect 487 -561 492 -521
rect 467 -567 472 -563
rect 478 -568 483 -566
rect 487 -568 492 -566
rect 511 -545 516 -539
rect 511 -557 516 -551
rect 511 -567 516 -563
rect 520 -533 525 -521
rect 520 -545 525 -539
rect 520 -557 525 -551
rect 540 -561 545 -521
rect 520 -567 525 -563
rect 531 -568 536 -566
rect 540 -568 545 -566
rect 564 -545 569 -539
rect 564 -557 569 -551
rect 564 -567 569 -563
rect 573 -533 578 -521
rect 573 -545 578 -539
rect 573 -557 578 -551
rect 593 -561 598 -521
rect 573 -567 578 -563
rect 584 -568 589 -566
rect 593 -568 598 -566
rect 617 -545 622 -539
rect 617 -557 622 -551
rect 617 -567 622 -563
rect 626 -533 631 -521
rect 626 -545 631 -539
rect 626 -557 631 -551
rect 646 -561 651 -521
rect 626 -567 631 -563
rect 637 -568 642 -566
rect 646 -568 651 -566
rect 670 -545 675 -539
rect 670 -557 675 -551
rect 670 -567 675 -563
rect 679 -533 684 -521
rect 679 -545 684 -539
rect 679 -557 684 -551
rect 699 -561 704 -521
rect 679 -567 684 -563
rect 690 -568 695 -566
rect 699 -568 704 -566
rect 723 -545 728 -539
rect 723 -557 728 -551
rect 723 -567 728 -563
rect 732 -533 737 -521
rect 732 -545 737 -539
rect 732 -557 737 -551
rect 752 -561 757 -521
rect 767 -521 772 -504
rect 732 -567 737 -563
rect 743 -568 748 -566
rect 752 -568 757 -566
rect 266 -586 271 -573
rect 276 -579 280 -573
rect 319 -586 324 -573
rect 329 -579 333 -573
rect 372 -586 377 -573
rect 382 -579 386 -573
rect 425 -586 430 -573
rect 435 -579 439 -573
rect 478 -586 483 -573
rect 488 -579 492 -573
rect 531 -586 536 -573
rect 541 -579 545 -573
rect 584 -586 589 -573
rect 594 -579 598 -573
rect 637 -586 642 -573
rect 647 -579 651 -573
rect 690 -586 695 -573
rect 700 -579 704 -573
rect 743 -586 748 -573
rect 753 -579 757 -573
rect -459 -599 -450 -593
rect -237 -594 -181 -593
rect -237 -598 -225 -594
rect -221 -598 -209 -594
rect -205 -598 -181 -594
rect -237 -599 -181 -598
rect 88 -587 767 -586
rect 88 -593 240 -587
rect 244 -593 250 -587
rect 254 -593 259 -587
rect 263 -593 267 -587
rect 271 -593 275 -587
rect 279 -593 283 -587
rect 287 -593 293 -587
rect 297 -593 303 -587
rect 307 -593 312 -587
rect 316 -593 320 -587
rect 324 -593 328 -587
rect 332 -593 336 -587
rect 340 -593 346 -587
rect 350 -593 356 -587
rect 360 -593 365 -587
rect 369 -593 373 -587
rect 377 -593 381 -587
rect 385 -593 389 -587
rect 393 -593 399 -587
rect 403 -593 409 -587
rect 413 -593 418 -587
rect 422 -593 426 -587
rect 430 -593 434 -587
rect 438 -593 442 -587
rect 446 -593 452 -587
rect 456 -593 462 -587
rect 466 -593 471 -587
rect 475 -593 479 -587
rect 483 -593 487 -587
rect 491 -593 495 -587
rect 499 -593 505 -587
rect 509 -593 515 -587
rect 519 -593 524 -587
rect 528 -593 532 -587
rect 536 -593 540 -587
rect 544 -593 548 -587
rect 552 -593 558 -587
rect 562 -593 568 -587
rect 572 -593 577 -587
rect 581 -593 585 -587
rect 589 -593 593 -587
rect 597 -593 601 -587
rect 605 -593 611 -587
rect 615 -593 621 -587
rect 625 -593 630 -587
rect 634 -593 638 -587
rect 642 -593 646 -587
rect 650 -593 654 -587
rect 658 -593 664 -587
rect 668 -593 674 -587
rect 678 -593 683 -587
rect 687 -593 691 -587
rect 695 -593 699 -587
rect 703 -593 707 -587
rect 711 -593 717 -587
rect 721 -593 727 -587
rect 731 -593 736 -587
rect 740 -593 744 -587
rect 748 -593 752 -587
rect 756 -593 760 -587
rect 764 -593 767 -587
rect 88 -594 767 -593
rect 88 -602 94 -594
rect -13 -606 24 -602
rect 28 -606 32 -602
rect 36 -606 40 -602
rect 44 -606 48 -602
rect 52 -606 56 -602
rect 60 -606 64 -602
rect 68 -606 72 -602
rect 76 -606 80 -602
rect 84 -606 88 -602
rect 92 -606 94 -602
rect 104 -606 105 -602
rect 109 -606 113 -602
rect 117 -606 121 -602
rect 125 -606 130 -602
rect 134 -606 138 -602
rect 142 -606 144 -602
rect -13 -611 -1 -606
rect -144 -620 -96 -619
rect -144 -626 -140 -620
rect -136 -626 -132 -620
rect -128 -626 -124 -620
rect -120 -626 -116 -620
rect -112 -626 -108 -620
rect -104 -626 -96 -620
rect -144 -627 -96 -626
rect -139 -632 -134 -627
rect -156 -648 -148 -642
rect -158 -656 -148 -651
rect -130 -657 -125 -642
rect -139 -665 -134 -662
rect -139 -672 -134 -670
rect -139 -690 -134 -677
rect -130 -665 -125 -662
rect -130 -672 -125 -670
rect -130 -683 -125 -677
rect -121 -657 -116 -642
rect -121 -665 -116 -662
rect -121 -672 -116 -670
rect -112 -657 -107 -648
rect -112 -665 -107 -662
rect 24 -651 28 -606
rect 24 -656 28 -655
rect 24 -661 28 -660
rect 24 -666 28 -665
rect 36 -655 40 -654
rect 36 -660 40 -659
rect 36 -665 40 -664
rect -112 -672 -107 -670
rect 36 -675 40 -669
rect 45 -651 49 -606
rect 73 -611 77 -606
rect 73 -616 77 -615
rect 73 -621 77 -620
rect 73 -626 77 -625
rect 73 -631 77 -630
rect 73 -636 77 -635
rect 73 -641 77 -640
rect 73 -646 77 -645
rect 45 -656 49 -655
rect 45 -661 49 -660
rect 45 -666 49 -665
rect 57 -655 61 -654
rect 57 -660 61 -659
rect 57 -665 61 -664
rect -121 -683 -116 -677
rect 35 -679 50 -675
rect -121 -687 -79 -683
rect -145 -691 -97 -690
rect -145 -697 -138 -691
rect -134 -697 -130 -691
rect -126 -697 -120 -691
rect -116 -697 -112 -691
rect -108 -697 -104 -691
rect -100 -697 -97 -691
rect -145 -698 -97 -697
rect 24 -697 28 -696
rect 24 -702 28 -701
rect 24 -707 28 -706
rect 16 -711 24 -708
rect 16 -712 28 -711
rect 36 -693 40 -679
rect 57 -680 61 -669
rect 73 -651 77 -650
rect 73 -656 77 -655
rect 73 -661 77 -660
rect 73 -666 77 -665
rect 85 -615 89 -614
rect 85 -620 89 -619
rect 85 -625 89 -624
rect 85 -630 89 -629
rect 85 -635 89 -634
rect 85 -640 89 -639
rect 85 -645 89 -644
rect 85 -650 89 -649
rect 85 -655 89 -654
rect 85 -660 89 -659
rect 85 -665 89 -664
rect 110 -653 114 -606
rect 110 -658 114 -657
rect 110 -663 114 -662
rect 89 -669 94 -665
rect 48 -687 50 -683
rect 82 -680 86 -678
rect 36 -698 40 -697
rect 36 -703 40 -702
rect 36 -708 40 -707
rect 45 -697 49 -696
rect 45 -702 49 -701
rect 45 -707 49 -706
rect 16 -727 20 -712
rect 35 -721 37 -717
rect 45 -727 49 -711
rect 57 -693 61 -684
rect 90 -689 94 -669
rect 110 -668 114 -667
rect 122 -657 126 -656
rect 122 -662 126 -661
rect 122 -667 126 -666
rect 122 -689 126 -671
rect 131 -653 135 -606
rect 131 -658 135 -657
rect 131 -663 135 -662
rect 131 -668 135 -667
rect 143 -652 147 -613
rect 312 -626 316 -619
rect 392 -627 396 -620
rect 472 -627 476 -616
rect 552 -627 556 -620
rect 632 -627 636 -620
rect 143 -657 147 -656
rect 143 -662 147 -661
rect 143 -667 147 -666
rect 57 -698 61 -697
rect 57 -703 61 -702
rect 57 -708 61 -707
rect 73 -693 113 -689
rect 122 -693 134 -689
rect 16 -731 52 -727
rect -13 -758 -1 -753
rect 20 -748 47 -744
rect 51 -748 66 -744
rect 20 -758 24 -748
rect -13 -762 15 -758
rect 19 -762 24 -758
rect 8 -770 12 -769
rect 8 -775 12 -774
rect 8 -780 12 -779
rect 8 -789 12 -784
rect 20 -766 24 -762
rect 20 -771 24 -770
rect 20 -776 24 -775
rect 20 -781 24 -780
rect 40 -764 44 -763
rect 40 -769 44 -768
rect 40 -774 44 -773
rect 40 -789 44 -778
rect 52 -760 56 -758
rect 52 -765 56 -764
rect 52 -770 56 -769
rect 52 -775 56 -774
rect 61 -764 65 -763
rect 61 -769 65 -768
rect 61 -774 65 -773
rect -2 -793 1 -789
rect 5 -793 9 -789
rect 13 -793 17 -789
rect 21 -793 25 -789
rect 29 -793 33 -789
rect 37 -793 41 -789
rect 45 -793 49 -789
rect 53 -793 57 -789
rect 61 -793 65 -778
rect 73 -760 77 -693
rect 73 -765 77 -764
rect 73 -770 77 -769
rect 73 -775 77 -774
rect 110 -702 114 -701
rect 110 -789 114 -706
rect 122 -698 126 -693
rect 122 -703 126 -702
rect 131 -702 135 -701
rect 131 -789 135 -706
rect 143 -698 147 -671
rect 143 -703 147 -702
rect 332 -633 348 -627
rect 360 -633 368 -627
rect 412 -633 428 -627
rect 440 -633 448 -627
rect 492 -633 508 -627
rect 520 -633 528 -627
rect 572 -633 588 -627
rect 600 -633 608 -627
rect 652 -633 668 -627
rect 680 -633 688 -627
rect 69 -793 73 -789
rect 77 -793 81 -789
rect 85 -793 87 -789
rect 100 -793 104 -789
rect 108 -793 112 -789
rect 116 -793 120 -789
rect 124 -793 129 -789
rect 133 -793 137 -789
rect 141 -793 145 -789
rect 149 -793 152 -789
rect 295 -811 299 -721
rect 312 -727 316 -716
rect 332 -727 336 -633
rect 352 -727 356 -717
rect 372 -811 376 -717
rect 392 -727 396 -717
rect 412 -727 416 -633
rect 432 -727 436 -717
rect 452 -811 456 -717
rect 472 -727 476 -717
rect 492 -727 496 -633
rect 512 -727 516 -717
rect 532 -811 536 -717
rect 552 -727 556 -717
rect 572 -727 576 -633
rect 592 -727 596 -717
rect 612 -811 616 -717
rect 632 -727 636 -717
rect 652 -727 656 -633
rect 672 -727 676 -717
rect 692 -722 696 -717
rect 295 -817 308 -811
rect 320 -817 328 -811
rect 372 -817 388 -811
rect 400 -817 408 -811
rect 452 -817 468 -811
rect 480 -817 488 -811
rect 532 -817 548 -811
rect 560 -817 568 -811
rect 612 -817 628 -811
rect 640 -817 648 -811
rect 352 -820 356 -817
rect 432 -820 436 -817
rect 512 -820 516 -817
rect 592 -820 596 -817
rect 672 -820 676 -817
<< m2contact >>
rect 1157 100 1161 106
rect -2 63 2 67
rect 228 63 232 67
rect 441 63 445 67
rect 669 63 673 67
rect 898 63 902 67
rect 236 50 240 54
rect 463 50 467 54
rect 685 50 689 54
rect 912 50 916 54
rect 449 40 453 44
rect 677 40 681 44
rect 905 40 909 44
rect -1 33 3 37
rect 221 36 225 40
rect 231 33 235 37
rect 456 33 460 37
rect 685 33 689 37
rect 918 33 922 37
rect 210 26 214 30
rect 441 9 445 13
rect 669 9 673 13
rect 898 7 902 11
rect 1132 0 1137 6
rect 1157 -27 1161 -21
rect -5 -77 -1 -73
rect 223 -77 227 -73
rect 451 -77 455 -73
rect 678 -77 682 -73
rect 907 -77 911 -73
rect 918 -73 922 -69
rect 1135 -78 1139 -73
rect 2 -87 6 -83
rect 1164 -87 1168 -83
rect -5 -94 -1 -90
rect 223 -94 227 -90
rect 451 -94 455 -90
rect 230 -98 234 -94
rect 678 -94 682 -90
rect -13 -102 -9 -98
rect 215 -102 219 -98
rect 443 -102 447 -98
rect 458 -99 462 -95
rect 914 -94 918 -90
rect 1135 -94 1139 -90
rect 686 -99 690 -95
rect 671 -103 675 -99
rect 899 -103 903 -99
rect 1127 -103 1131 -99
rect 1149 -127 1153 -121
rect 1157 -153 1161 -147
rect 918 -183 922 -179
rect 2 -190 6 -186
rect 230 -190 234 -186
rect 458 -190 462 -186
rect 686 -190 690 -186
rect 4 -203 8 -199
rect 6 -213 10 -209
rect 233 -203 237 -199
rect 234 -213 238 -209
rect 228 -220 232 -216
rect 461 -203 465 -199
rect 462 -213 466 -209
rect 456 -220 460 -216
rect 688 -203 692 -199
rect 690 -213 694 -209
rect 684 -220 688 -216
rect 916 -203 920 -199
rect 918 -213 922 -209
rect 912 -220 916 -216
rect 1132 -253 1137 -247
rect 1134 -273 1138 -267
rect 221 -302 225 -298
rect 449 -303 453 -299
rect 677 -303 681 -299
rect 905 -303 909 -299
rect 1134 -310 1138 -306
rect 466 -319 470 -315
rect 693 -319 697 -315
rect 920 -319 924 -315
rect -237 -331 -233 -327
rect -449 -340 -445 -336
rect -11 -331 -7 -327
rect -222 -340 -218 -336
rect 222 -323 226 -319
rect 221 -333 225 -329
rect 451 -323 455 -319
rect 448 -333 452 -329
rect 676 -323 680 -319
rect 676 -333 680 -329
rect 906 -323 910 -319
rect 905 -333 909 -329
rect 1133 -323 1137 -319
rect 1140 -333 1144 -329
rect 237 -340 241 -336
rect 1 -351 5 -346
rect 1133 -361 1137 -357
rect 1155 -373 1159 -367
rect -241 -436 -237 -432
rect -453 -444 -449 -440
rect -242 -453 -238 -449
rect -440 -477 -436 -473
rect -227 -432 -223 -428
rect 1 -391 5 -386
rect 565 -393 569 -389
rect 959 -393 963 -389
rect 1163 -393 1167 -389
rect -227 -444 -223 -440
rect -15 -453 -11 -449
rect 1155 -408 1159 -404
rect 480 -414 484 -410
rect 321 -465 325 -461
rect -210 -543 -206 -541
rect -210 -545 -206 -543
rect -446 -549 -442 -545
rect -240 -557 -236 -553
rect -230 -559 -226 -555
rect -452 -566 -448 -562
rect -196 -570 -192 -566
rect 374 -465 378 -461
rect 427 -466 431 -461
rect 1155 -415 1159 -411
rect 1155 -422 1159 -418
rect 1155 -429 1159 -425
rect 1155 -436 1159 -432
rect 1155 -443 1159 -439
rect 1155 -450 1159 -446
rect 586 -455 590 -451
rect 533 -467 537 -463
rect 1155 -457 1159 -453
rect 1155 -464 1159 -460
rect 639 -474 643 -470
rect 692 -471 696 -466
rect 745 -478 749 -473
rect 231 -533 236 -527
rect 246 -533 251 -527
rect 255 -573 260 -567
rect 299 -533 304 -527
rect 308 -573 313 -567
rect 352 -533 357 -527
rect 361 -573 366 -567
rect 405 -533 410 -527
rect 414 -573 419 -567
rect 458 -533 463 -527
rect 467 -573 472 -567
rect 511 -533 516 -527
rect 520 -573 525 -567
rect 564 -533 569 -527
rect 573 -573 578 -567
rect 617 -533 622 -527
rect 626 -573 631 -567
rect 670 -533 675 -527
rect 679 -573 684 -567
rect 723 -533 728 -527
rect 767 -527 772 -521
rect 732 -573 737 -567
rect -148 -648 -143 -642
rect -162 -656 -158 -651
rect -112 -648 -107 -642
rect -79 -687 -75 -683
rect 44 -687 48 -683
rect 57 -684 61 -680
rect 82 -684 86 -680
rect 37 -721 41 -717
rect 143 -613 147 -609
rect 312 -619 316 -615
rect 392 -620 396 -616
rect 467 -620 472 -616
rect 552 -620 556 -616
rect 632 -620 636 -616
rect 52 -731 56 -727
rect 52 -758 56 -754
rect 295 -721 299 -717
rect 692 -727 696 -722
rect 352 -824 356 -820
rect 432 -824 436 -820
rect 512 -824 516 -820
rect 592 -824 596 -820
rect 672 -824 676 -820
<< metal2 >>
rect -10 63 -2 67
rect 2 63 7 67
rect 210 63 228 67
rect -1 -3 3 33
rect 210 30 214 63
rect 233 50 236 54
rect 221 31 225 36
rect 231 -3 235 33
rect 441 13 445 63
rect 460 50 463 54
rect 449 33 453 40
rect 456 -3 460 33
rect 669 13 673 63
rect 685 45 689 50
rect 677 35 681 40
rect 685 -3 689 33
rect 898 11 902 63
rect 912 44 916 50
rect 905 34 909 40
rect 898 6 902 7
rect 918 -3 922 33
rect 1137 0 1153 6
rect -253 -7 1146 -3
rect -253 -254 -249 -7
rect -13 -64 -9 -60
rect -5 -83 -1 -77
rect 223 -83 227 -77
rect 451 -83 455 -77
rect 678 -83 682 -77
rect 907 -83 911 -77
rect 918 -77 922 -73
rect 1135 -82 1139 -78
rect -18 -102 -13 -98
rect -5 -130 -1 -94
rect 2 -91 6 -87
rect 2 -103 6 -95
rect 210 -102 215 -98
rect 223 -130 227 -94
rect 230 -102 234 -98
rect 438 -102 443 -98
rect 230 -114 234 -106
rect 451 -130 455 -94
rect 458 -103 462 -99
rect 666 -103 671 -99
rect 458 -115 462 -107
rect 678 -130 682 -94
rect 686 -103 690 -99
rect 894 -103 899 -99
rect 686 -115 690 -107
rect 914 -130 918 -94
rect 1122 -103 1127 -99
rect 1135 -130 1139 -94
rect 1142 -130 1146 -7
rect -5 -134 1146 -130
rect 1149 -121 1153 0
rect 686 -167 690 -166
rect 230 -178 234 -177
rect 2 -186 6 -182
rect 230 -186 234 -182
rect 458 -186 462 -173
rect 686 -186 690 -171
rect 918 -179 922 -166
rect -4 -203 4 -199
rect 219 -203 233 -199
rect 447 -203 461 -199
rect 676 -203 688 -199
rect 903 -203 916 -199
rect -4 -232 0 -203
rect -450 -258 -249 -254
rect 6 -257 10 -213
rect 219 -233 223 -203
rect 228 -224 232 -220
rect 235 -257 238 -213
rect 447 -225 451 -203
rect 456 -223 460 -220
rect 463 -257 466 -213
rect 676 -224 680 -203
rect 684 -222 688 -220
rect 691 -257 694 -213
rect 903 -230 907 -203
rect 912 -221 916 -220
rect 919 -257 922 -213
rect 1149 -247 1153 -127
rect 1157 -21 1161 100
rect 1157 -147 1161 -27
rect 1164 -94 1168 -87
rect 1157 -196 1161 -153
rect 1137 -253 1159 -247
rect -450 -336 -446 -258
rect 6 -261 1152 -257
rect 1138 -273 1141 -269
rect 221 -298 225 -294
rect 449 -299 453 -296
rect 677 -299 681 -295
rect 905 -299 909 -295
rect 1138 -310 1141 -306
rect 226 -323 234 -319
rect 455 -323 462 -319
rect -245 -331 -237 -329
rect -245 -333 -233 -331
rect -19 -331 -11 -329
rect -19 -333 -7 -331
rect -237 -336 -233 -333
rect -450 -340 -449 -336
rect -237 -340 -222 -336
rect -234 -432 -227 -428
rect -241 -442 -237 -436
rect -449 -444 -441 -442
rect -453 -446 -441 -444
rect -453 -562 -449 -446
rect -234 -449 -230 -432
rect -223 -444 -215 -442
rect -227 -446 -215 -444
rect -14 -449 -10 -333
rect 1 -386 5 -351
rect 221 -376 225 -333
rect 230 -354 234 -323
rect 237 -342 241 -340
rect 448 -376 452 -333
rect 458 -349 462 -323
rect 466 -321 470 -319
rect 680 -323 690 -319
rect 676 -376 680 -333
rect 686 -348 690 -323
rect 693 -320 697 -319
rect 910 -323 916 -319
rect 912 -325 916 -323
rect 920 -320 924 -319
rect 905 -376 909 -333
rect 1133 -357 1137 -323
rect 1148 -329 1152 -261
rect 1144 -333 1152 -329
rect 1148 -376 1152 -333
rect 1155 -367 1159 -253
rect 13 -380 1152 -376
rect -238 -453 -230 -449
rect -11 -453 -10 -449
rect -440 -486 -436 -477
rect -440 -490 -226 -486
rect -446 -543 -430 -539
rect -446 -545 -442 -543
rect -248 -557 -240 -555
rect -248 -559 -236 -557
rect -230 -555 -226 -490
rect -206 -545 -158 -541
rect -453 -566 -452 -562
rect -239 -570 -196 -566
rect -162 -651 -158 -545
rect 13 -580 17 -380
rect 561 -393 565 -389
rect 963 -393 1144 -389
rect 1148 -393 1163 -389
rect 950 -410 954 -394
rect 1130 -404 1134 -401
rect 1130 -408 1155 -404
rect 484 -414 954 -410
rect 950 -425 954 -414
rect 1130 -415 1155 -411
rect 1130 -422 1155 -418
rect 950 -429 1155 -425
rect 1148 -436 1155 -432
rect 321 -439 325 -438
rect 1148 -443 1155 -439
rect 321 -461 325 -443
rect 374 -461 378 -447
rect 427 -461 431 -448
rect 586 -451 590 -443
rect 1148 -450 1155 -446
rect 533 -463 537 -456
rect 639 -470 643 -458
rect 1148 -457 1155 -453
rect 692 -466 696 -460
rect 1148 -464 1155 -460
rect 745 -473 749 -467
rect 236 -533 246 -527
rect 251 -533 299 -527
rect 304 -533 352 -527
rect 357 -533 405 -527
rect 410 -533 458 -527
rect 463 -533 511 -527
rect 516 -533 564 -527
rect 569 -533 617 -527
rect 622 -533 670 -527
rect 675 -533 723 -527
rect 728 -533 756 -527
rect 13 -584 147 -580
rect 143 -609 147 -584
rect 255 -615 260 -573
rect 308 -605 313 -573
rect 308 -610 356 -605
rect 255 -619 312 -615
rect -143 -648 -112 -642
rect -75 -687 44 -683
rect 61 -684 82 -680
rect 41 -721 295 -717
rect 52 -754 56 -731
rect 352 -820 356 -610
rect 361 -616 366 -573
rect 414 -611 419 -573
rect 414 -616 436 -611
rect 361 -620 392 -616
rect 432 -820 436 -616
rect 467 -616 472 -573
rect 520 -616 525 -573
rect 573 -616 578 -573
rect 626 -605 631 -573
rect 679 -602 684 -573
rect 512 -620 525 -616
rect 556 -620 578 -616
rect 592 -610 631 -605
rect 646 -606 684 -602
rect 512 -820 516 -620
rect 592 -820 596 -610
rect 646 -616 650 -606
rect 636 -620 650 -616
rect 732 -617 737 -573
rect 672 -621 737 -617
rect 672 -820 676 -621
rect 767 -722 772 -527
rect 696 -727 772 -722
<< m3contact >>
rect -14 62 -10 67
rect 229 50 233 54
rect 221 27 225 31
rect 456 50 460 54
rect 449 29 453 33
rect 685 41 689 45
rect 677 31 681 35
rect 912 40 916 44
rect 905 30 909 34
rect -22 -64 -18 -60
rect 206 -64 210 -60
rect 434 -64 438 -60
rect 662 -64 666 -60
rect 890 -64 894 -60
rect 1118 -64 1122 -60
rect -5 -87 -1 -83
rect 223 -87 227 -83
rect 451 -87 455 -83
rect 678 -87 682 -83
rect 918 -81 922 -77
rect 907 -87 911 -83
rect 1135 -87 1139 -82
rect -22 -102 -18 -98
rect 2 -95 6 -91
rect 206 -102 210 -98
rect 434 -102 438 -98
rect 230 -106 234 -102
rect 662 -103 666 -99
rect 458 -107 462 -103
rect 890 -103 894 -99
rect 686 -107 690 -103
rect 1118 -103 1122 -99
rect 918 -166 922 -162
rect 458 -173 462 -169
rect 2 -182 6 -178
rect 230 -182 234 -178
rect 686 -171 690 -167
rect -4 -236 0 -232
rect 228 -228 232 -224
rect 219 -237 223 -233
rect 447 -229 451 -225
rect 456 -227 460 -223
rect 676 -228 680 -224
rect 684 -226 688 -222
rect 912 -225 916 -221
rect 903 -234 907 -230
rect 1164 -98 1168 -94
rect 1157 -200 1161 -196
rect 1141 -273 1145 -269
rect 221 -294 225 -290
rect 449 -296 453 -292
rect 677 -295 681 -291
rect 905 -295 909 -291
rect 1141 -310 1145 -306
rect -249 -333 -245 -329
rect -23 -333 -19 -329
rect -441 -446 -437 -442
rect -241 -446 -237 -442
rect -215 -446 -211 -442
rect 237 -346 241 -342
rect 230 -358 234 -354
rect 466 -325 470 -321
rect 458 -353 462 -349
rect 693 -324 697 -320
rect 920 -324 924 -320
rect 912 -329 916 -325
rect 686 -352 690 -348
rect -430 -543 -426 -539
rect -252 -559 -248 -555
rect -243 -570 -239 -566
rect 557 -393 561 -389
rect 950 -394 954 -389
rect 1144 -393 1148 -389
rect 1130 -401 1134 -397
rect 1126 -415 1130 -411
rect 1126 -422 1130 -418
rect 1144 -436 1148 -432
rect 321 -443 325 -439
rect 586 -443 590 -439
rect 1144 -443 1148 -439
rect 374 -447 378 -443
rect 427 -448 431 -443
rect 1144 -450 1148 -446
rect 533 -456 537 -452
rect 639 -458 643 -454
rect 692 -460 696 -455
rect 1144 -457 1148 -453
rect 745 -467 749 -462
rect 1144 -464 1148 -460
<< metal3 >>
rect -14 -10 -10 62
rect 221 20 225 27
rect 229 -10 233 50
rect 449 25 453 29
rect 456 -10 460 50
rect 677 27 681 31
rect 685 -10 689 41
rect 905 26 909 30
rect 912 -10 916 40
rect -14 -14 1159 -10
rect -22 -98 -18 -64
rect -5 -137 -1 -87
rect 2 -99 6 -95
rect 206 -98 210 -64
rect 223 -137 227 -87
rect 434 -98 438 -64
rect 230 -110 234 -106
rect 451 -137 455 -87
rect 662 -99 666 -64
rect 458 -111 462 -107
rect 678 -137 682 -87
rect 890 -99 894 -64
rect 686 -111 690 -107
rect 907 -137 911 -87
rect 918 -86 922 -81
rect 1118 -99 1122 -64
rect 1135 -137 1139 -87
rect 1155 -137 1159 -14
rect 1164 -103 1168 -98
rect -230 -141 1159 -137
rect -230 -260 -226 -141
rect 2 -178 6 -165
rect 230 -178 234 -162
rect 458 -169 462 -164
rect 686 -167 690 -162
rect 918 -162 922 -158
rect 1157 -205 1161 -200
rect 228 -230 232 -228
rect -4 -260 0 -236
rect 219 -260 223 -237
rect 447 -260 451 -229
rect 456 -229 460 -227
rect 676 -260 680 -228
rect 684 -228 688 -226
rect 912 -228 916 -225
rect 903 -260 907 -234
rect -230 -264 1177 -260
rect 1145 -273 1150 -269
rect 221 -290 225 -284
rect 449 -292 453 -285
rect 677 -291 681 -287
rect 905 -291 909 -284
rect 1145 -310 1164 -306
rect -346 -333 -249 -329
rect -120 -333 -23 -329
rect 466 -332 470 -325
rect 693 -333 697 -324
rect 237 -349 241 -346
rect 230 -382 234 -358
rect 458 -382 462 -353
rect 686 -382 690 -352
rect 912 -382 916 -329
rect 920 -335 924 -324
rect 1173 -382 1177 -264
rect 230 -386 1177 -382
rect 548 -393 557 -389
rect 924 -394 950 -389
rect 237 -397 241 -394
rect 237 -401 1130 -397
rect 321 -439 325 -401
rect -437 -446 -340 -442
rect -243 -446 -241 -442
rect -211 -446 -114 -442
rect 374 -443 378 -411
rect -243 -539 -239 -446
rect 1110 -415 1126 -411
rect 427 -443 431 -415
rect 1106 -422 1126 -418
rect 1144 -432 1148 -393
rect 590 -443 1052 -439
rect 1056 -443 1144 -439
rect 533 -452 537 -447
rect 639 -454 643 -450
rect 1042 -450 1144 -446
rect 692 -455 696 -451
rect 745 -462 749 -455
rect 1032 -457 1144 -453
rect 1017 -464 1144 -460
rect -426 -543 -239 -539
rect -349 -559 -252 -555
rect -243 -566 -239 -543
<< m4contact >>
rect 221 16 225 20
rect 449 21 453 25
rect 677 23 681 27
rect 905 22 909 26
rect 2 -103 6 -99
rect 230 -114 234 -110
rect 458 -115 462 -111
rect 686 -115 690 -111
rect 918 -90 922 -86
rect 1164 -107 1168 -103
rect 918 -158 922 -154
rect 2 -165 6 -161
rect 230 -162 234 -158
rect 458 -164 462 -160
rect 686 -162 690 -158
rect 1157 -209 1161 -205
rect 228 -234 232 -230
rect 456 -233 460 -229
rect 684 -232 688 -228
rect 912 -232 916 -228
rect 1150 -273 1154 -269
rect 221 -284 225 -280
rect 449 -285 453 -281
rect 677 -287 681 -283
rect 905 -284 909 -280
rect 1164 -310 1168 -306
rect 466 -336 470 -332
rect 693 -337 697 -333
rect 237 -353 241 -349
rect 920 -339 924 -335
rect 237 -394 241 -389
rect 544 -393 548 -389
rect 920 -394 924 -389
rect 374 -411 378 -407
rect 1110 -411 1114 -407
rect 427 -415 431 -411
rect 1102 -422 1106 -418
rect 1052 -443 1056 -439
rect 533 -447 537 -443
rect 639 -450 643 -446
rect 692 -451 696 -446
rect 1038 -450 1042 -446
rect 745 -455 749 -451
rect 1028 -457 1032 -453
rect 1013 -464 1017 -460
<< metal4 >>
rect 2 -161 6 -103
rect 221 -280 225 16
rect 230 -158 234 -114
rect 228 -236 232 -234
rect 449 -281 453 21
rect 458 -160 462 -115
rect 456 -236 460 -233
rect 677 -283 681 23
rect 686 -158 690 -115
rect 684 -234 688 -232
rect 905 -280 909 22
rect 918 -154 922 -90
rect 912 -235 916 -232
rect 1157 -269 1161 -209
rect 1154 -273 1161 -269
rect 1164 -306 1168 -107
rect 237 -389 241 -353
rect 466 -403 470 -336
rect 693 -383 697 -337
rect 920 -389 924 -339
rect 537 -393 544 -389
rect 374 -407 1114 -403
rect 431 -415 693 -411
rect 533 -443 537 -422
rect 639 -429 684 -425
rect 639 -446 643 -429
rect 692 -446 696 -436
rect 745 -451 749 -443
rect 1013 -460 1017 -443
rect 1028 -453 1032 -436
rect 1038 -446 1042 -429
rect 1052 -439 1056 -415
rect 1092 -422 1102 -418
<< m5contact >>
rect 228 -240 232 -236
rect 456 -240 460 -236
rect 684 -238 688 -234
rect 912 -239 916 -235
rect 693 -388 697 -383
rect 533 -393 537 -389
rect 693 -415 697 -411
rect 1052 -415 1056 -411
rect 533 -422 537 -418
rect 684 -429 688 -425
rect 1038 -429 1042 -425
rect 692 -436 696 -432
rect 1028 -436 1032 -432
rect 745 -443 749 -439
rect 1013 -443 1017 -439
rect 1088 -422 1092 -418
<< metal5 >>
rect 228 -439 232 -240
rect 456 -432 460 -240
rect 533 -418 537 -393
rect 684 -425 688 -238
rect 693 -411 697 -388
rect 912 -386 916 -239
rect 912 -390 1056 -386
rect 1052 -411 1056 -390
rect 693 -418 697 -415
rect 693 -422 1088 -418
rect 688 -429 1038 -425
rect 456 -436 692 -432
rect 696 -436 1028 -432
rect 228 -443 745 -439
rect 749 -443 1013 -439
<< pseudo_rnwell >>
rect -14 -611 0 -610
rect -14 -753 -13 -611
rect -1 -753 0 -611
rect 307 -626 321 -625
rect 307 -716 308 -626
rect 320 -716 321 -626
rect 307 -717 321 -716
rect 347 -627 361 -626
rect 347 -717 348 -627
rect 360 -717 361 -627
rect 347 -718 361 -717
rect 367 -627 381 -626
rect 367 -717 368 -627
rect 380 -717 381 -627
rect 367 -718 381 -717
rect 387 -627 401 -626
rect 387 -717 388 -627
rect 400 -717 401 -627
rect 387 -718 401 -717
rect 427 -627 441 -626
rect 427 -717 428 -627
rect 440 -717 441 -627
rect 427 -718 441 -717
rect 447 -627 461 -626
rect 447 -717 448 -627
rect 460 -717 461 -627
rect 447 -718 461 -717
rect 467 -627 481 -626
rect 467 -717 468 -627
rect 480 -717 481 -627
rect 467 -718 481 -717
rect 507 -627 521 -626
rect 507 -717 508 -627
rect 520 -717 521 -627
rect 507 -718 521 -717
rect 527 -627 541 -626
rect 527 -717 528 -627
rect 540 -717 541 -627
rect 527 -718 541 -717
rect 547 -627 561 -626
rect 547 -717 548 -627
rect 560 -717 561 -627
rect 547 -718 561 -717
rect 587 -627 601 -626
rect 587 -717 588 -627
rect 600 -717 601 -627
rect 587 -718 601 -717
rect 607 -627 621 -626
rect 607 -717 608 -627
rect 620 -717 621 -627
rect 607 -718 621 -717
rect 627 -627 641 -626
rect 627 -717 628 -627
rect 640 -717 641 -627
rect 627 -718 641 -717
rect 667 -627 681 -626
rect 667 -717 668 -627
rect 680 -717 681 -627
rect 667 -718 681 -717
rect 687 -627 701 -626
rect 687 -717 688 -627
rect 700 -717 701 -627
rect 687 -718 701 -717
rect 307 -727 321 -726
rect -14 -754 0 -753
rect 307 -817 308 -727
rect 320 -817 321 -727
rect 307 -818 321 -817
rect 327 -727 341 -726
rect 327 -817 328 -727
rect 340 -817 341 -727
rect 327 -818 341 -817
rect 347 -727 361 -726
rect 347 -817 348 -727
rect 360 -817 361 -727
rect 347 -818 361 -817
rect 387 -727 401 -726
rect 387 -817 388 -727
rect 400 -817 401 -727
rect 387 -818 401 -817
rect 407 -727 421 -726
rect 407 -817 408 -727
rect 420 -817 421 -727
rect 407 -818 421 -817
rect 427 -727 441 -726
rect 427 -817 428 -727
rect 440 -817 441 -727
rect 427 -818 441 -817
rect 467 -727 481 -726
rect 467 -817 468 -727
rect 480 -817 481 -727
rect 467 -818 481 -817
rect 487 -727 501 -726
rect 487 -817 488 -727
rect 500 -817 501 -727
rect 487 -818 501 -817
rect 507 -727 521 -726
rect 507 -817 508 -727
rect 520 -817 521 -727
rect 507 -818 521 -817
rect 547 -727 561 -726
rect 547 -817 548 -727
rect 560 -817 561 -727
rect 547 -818 561 -817
rect 567 -727 581 -726
rect 567 -817 568 -727
rect 580 -817 581 -727
rect 567 -818 581 -817
rect 587 -727 601 -726
rect 587 -817 588 -727
rect 600 -817 601 -727
rect 587 -818 601 -817
rect 627 -727 641 -726
rect 627 -817 628 -727
rect 640 -817 641 -727
rect 627 -818 641 -817
rect 647 -727 661 -726
rect 647 -817 648 -727
rect 660 -817 661 -727
rect 647 -818 661 -817
rect 667 -727 681 -726
rect 667 -817 668 -727
rect 680 -817 681 -727
rect 667 -818 681 -817
<< rnwell >>
rect -13 -747 -1 -617
rect 308 -710 320 -632
rect 348 -711 360 -633
rect 368 -711 380 -633
rect 388 -711 400 -633
rect 428 -711 440 -633
rect 448 -711 460 -633
rect 468 -711 480 -633
rect 508 -711 520 -633
rect 528 -711 540 -633
rect 548 -711 560 -633
rect 588 -711 600 -633
rect 608 -711 620 -633
rect 628 -711 640 -633
rect 668 -711 680 -633
rect 688 -711 700 -633
rect 308 -811 320 -733
rect 328 -811 340 -733
rect 348 -811 360 -733
rect 388 -811 400 -733
rect 408 -811 420 -733
rect 428 -811 440 -733
rect 468 -811 480 -733
rect 488 -811 500 -733
rect 508 -811 520 -733
rect 548 -811 560 -733
rect 568 -811 580 -733
rect 588 -811 600 -733
rect 628 -811 640 -733
rect 648 -811 660 -733
rect 668 -811 680 -733
use dffsr  dffsr_26
timestamp 1597999042
transform 1 0 -415 0 1 -596
box -38 -3 184 105
use dffsr  dffsr_25
timestamp 1597999042
transform -1 0 -274 0 1 -483
box -38 -3 184 105
use dffsr  dffsr_24
timestamp 1597999042
transform -1 0 -48 0 1 -483
box -38 -3 184 105
use dffsr  dffsr_22
timestamp 1597999042
transform 1 0 -412 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_23
timestamp 1597999042
transform 1 0 -186 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_11
timestamp 1597999042
transform 1 0 -186 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_21
timestamp 1597999042
transform -1 0 188 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_12
timestamp 1597999042
transform 1 0 42 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_13
timestamp 1597999042
transform 1 0 270 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_20
timestamp 1597999042
transform -1 0 416 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_14
timestamp 1597999042
transform 1 0 498 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_19
timestamp 1597999042
transform -1 0 644 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_15
timestamp 1597999042
transform 1 0 726 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_18
timestamp 1597999042
transform -1 0 872 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_16
timestamp 1597999042
transform 1 0 954 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_17
timestamp 1597999042
transform -1 0 1100 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_10
timestamp 1597999042
transform -1 0 -40 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_9
timestamp 1597999042
transform -1 0 188 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_0
timestamp 1597999042
transform 1 0 38 0 1 3
box -38 -3 184 105
use dffsr  dffsr_8
timestamp 1597999042
transform -1 0 416 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_1
timestamp 1597999042
transform 1 0 267 0 1 3
box -38 -3 184 105
use dffsr  dffsr_7
timestamp 1597999042
transform -1 0 644 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_2
timestamp 1597999042
transform 1 0 495 0 1 3
box -38 -3 184 105
use dffsr  dffsr_6
timestamp 1597999042
transform -1 0 872 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_3
timestamp 1597999042
transform 1 0 723 0 1 3
box -38 -3 184 105
use dffsr  dffsr_5
timestamp 1597999042
transform -1 0 1100 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_4
timestamp 1597999042
transform 1 0 954 0 1 3
box -38 -3 184 105
<< labels >>
rlabel metal2 428 -6 428 -6 1 CLK
rlabel metal3 416 -12 416 -12 1 SOC
rlabel metal1 912 103 912 103 5 1
rlabel metal1 909 3 909 3 1 0
rlabel metal1 230 -85 230 -85 1 q9
rlabel metal1 908 54 908 54 1 q4
rlabel metal1 913 -85 913 -85 1 q6
rlabel metal1 684 -86 684 -86 1 q7
rlabel metal1 457 -85 457 -85 1 q8
rlabel metal1 0 -85 0 -85 1 q10
rlabel metal1 -227 -71 -227 -71 3 EOC
rlabel metal1 1148 56 1148 56 1 q5
rlabel metal1 452 56 452 56 1 q2
rlabel metal1 224 56 224 56 1 q1
rlabel metal1 227 -197 227 -197 1 D0
rlabel metal1 455 -197 455 -197 1 D1
rlabel metal1 683 -197 683 -197 1 D2
rlabel metal1 911 -198 911 -198 1 D3
rlabel metal1 680 56 680 56 1 q3
rlabel metal1 231 -317 231 -317 1 D8
rlabel metal1 459 -318 459 -318 1 D7
rlabel metal1 687 -317 687 -317 1 D6
rlabel metal1 915 -317 915 -317 1 D5
rlabel metal1 2 -317 2 -317 1 D9
rlabel metal1 228 -530 228 -530 3 vref
rlabel metal1 1145 -198 1145 -198 1 D4
rlabel metal1 247 -499 247 -499 1 0
rlabel metal1 248 -590 248 -590 1 vdda
rlabel metal2 223 -378 223 -378 1 comp
rlabel metal1 297 -814 297 -814 5 out_dac
rlabel metal1 120 -604 120 -604 1 1
rlabel metal1 19 -604 19 -604 1 vdda
rlabel metal1 -1 -791 -1 -791 1 0
rlabel metal1 -95 -685 -95 -685 7 out_sam
rlabel metal1 -125 -622 -125 -622 5 0
rlabel metal1 -150 -645 -150 -645 1 in
rlabel metal1 -132 -694 -132 -694 1 vdda
rlabel metal1 118 -790 118 -790 1 0
<< end >>
