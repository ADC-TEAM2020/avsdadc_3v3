* 10-Bit SAR ADC
.include osu018.lib
*****************************************
.subckt sample 1 0 in clk1 out
M1 in cbar out 1 pfet l=0.2u w=2u
M2 in clk1 out 0 nfet l=0.2u w=1u
M3 cbar clk1 1 1 pfet l=0.2u w=2u
M4 cbar clk1 0 0 nfet l=0.2u w=1u
C1 out 0 1p
.ends sample

.subckt AND N001 0 N003 N004 OUT
M1 N001 N003 N002 N001 pfet l=0.2u w=2u
M2 N001 N004 N002 N001 pfet l=0.2u w=2u
M3 N002 N003 N005 0 nfet l=0.2u w=1u
M5 N001 N002 OUT N001 pfet l=0.2u w=2u
M6 OUT N002 0 0 nfet l=0.2u w=1u
M4 N005 N004 0 0 nfet l=0.2u w=1u
.ends AND

*****clkDivider24*****

.subckt clkdivider N001 0 N008 Q4
XU1 0 N001 N003 0 0 Q0 N003 N008 DFFSR
XU2 0 N001 N004 0 0 Q1 N004 N003 DFFSR
XU3 0 N001 N005 0 0 Q2 N005 N004 DFFSR
XU4 0 N001 N006 0 N002 Q3 N006 Q2 DFFSR
XU5 0 N001 N007 0 N002 Q4 N007 N006 DFFSR
XU6 N001 0 Q3 Q4 N002 AND
.ends clkdivider


.subckt DFFSR 0 1 D S_ R_ Q Q_bar CLK
Msp S S_ 1 1 pfet w=2u l=0.2u
Msn S S_ 0 0 nfet w=1u l=0.2u
Mrp R R_ 1 1 pfet w=2u l=0.2u
Mrn R R_ 0 0 nfet w=1u l=0.2u
M0 a R 1 1 pfet w=2u l=0.2u
M1 1 b a 1 pfet w=2u l=0.2u
M2 b c 1 1 pfet w=2u l=0.2u
M3 1 S b 1 pfet w=2u l=0.2u
M4 c dd a 1 pfet w=1u l=0.2u
M5 e f c 1 pfet w=1u l=0.2u
M6 1 D e 1 pfet w=2u l=0.2u
M7 1 dd f 1 pfet w=2u l=0.2u
M8 dd CLK 1 1 pfet w=2u l=0.2u
M9 g dd b 1 pfet w=1u l=0.2u
M10 h f g 1 pfet w=1u l=0.2u
M11 Q_bar g 1 1 pfet w=2u l=0.2u
M12 1 R Q_bar 1 pfet w=2u l=0.2u
M13 h Q_bar 1 1 pfet w=2u l=0.2u
M14 1 S h 1 pfet w=2u l=0.2u
M15 1 Q_bar Q 1 pfet w=2u l=0.2u
M16 j R a 0 nfet w=2u l=0.2u
M17 0 b j 0 nfet w=2u l=0.2u
M18 k c 0 0 nfet w=2u l=0.2u
M19 b S k 0 nfet w=2u l=0.2u
M20 c f a 0 nfet w=1u l=0.2u
M21 e dd c 0 nfet w=1u l=0.2u
M22 0 D e 0 nfet w=1u l=0.2u
M23 0 dd f 0 nfet w=1u l=0.2u
M24 dd CLK 0 0 nfet w=1u l=0.2u
M25 g f b 0 nfet w=1u l=0.2u
M26 h dd g 0 nfet w=1u l=0.2u
M27 l g Q_bar 0 nfet w=2u l=0.2u
M28 0 R l 0 nfet w=2u l=0.2u
M29 m Q_bar 0 0 nfet w=2u l=0.2u
M30 h S m 0 nfet w=2u l=0.2u
M31 0 Q_bar Q 0 nfet w=1u l=0.2u
.ends DFFSR

***Comparator***
.subckt comparator N001 N002 0 N006 N005 Vout
M1 N001 N003 N003 N001 pfet l=180n w=240n m=1
M2 N001 N003 N004 N001 pfet l=200n w=240n m=1
M3 N003 N005 N008 0 nfet l=200n w=240n m=1
M4 N004 N006 N008 0 nfet l=200n w=240n m=1
M5 N001 N004 N009 N001 pfet l=200n w=240n m=1
M6 N009 N007 0 0 nfet l=200n w=240n m=1
M7 N008 N007 0 0 nfet l=200n w=240n m=1
M8 N002 N009 N010 N002 pfet l=200n w=240n
M9 N002 N010 Vout N002 pfet l=200n w=240n
M10 N010 N009 0 0 nfet l=200n w=240n
M11 Vout N010 0 0 nfet l=200n w=240n
R1 N001 N007 2MEG
M13 N007 N007 0 0 nfet l=0.2u w=2.5u
.ends comparator

***SAR Logic***

.subckt SAR VDD 0 RESET CLK COMP D9 D8 D7 D6 D5 D4 D3 D2 D1 D0 EOC
XU1 0 VDD 0 RESET 0 N001 q1 CLK DFFSR
XU2 0 VDD N001 0 RESET N002 q2 CLK DFFSR
XU3 0 VDD N002 0 RESET N003 q3 CLK DFFSR
XU4 0 VDD N003 0 RESET N004 q4 CLK DFFSR
XU5 0 VDD N004 0 RESET N005 q5 CLK DFFSR
XU6 0 VDD N005 0 RESET N006 q6 CLK DFFSR
XU7 0 VDD N006 0 RESET N007 q7 CLK DFFSR
XU8 0 VDD N007 0 RESET N008 q8 CLK DFFSR
XU9 0 VDD N008 0 RESET N009 q9 CLK DFFSR
XU10 0 VDD N009 0 RESET N010 q10 CLK DFFSR
XU11 0 VDD N010 0 RESET EOC q11 CLK DFFSR
XU12 0 VDD COMP N010 RESET D0 q12 N011 DFFSR
XU13 0 VDD COMP N009 RESET D1 q13 D0 DFFSR
XU14 0 VDD COMP N008 RESET D2 q14 D1 DFFSR
XU15 0 VDD COMP N007 RESET D3 q15 D2 DFFSR
XU16 0 VDD COMP N006 RESET D4 q16 D3 DFFSR
XU17 0 VDD COMP N005 RESET D5 q17 D4 DFFSR
XU18 0 VDD COMP N004 RESET D6 q18 D5 DFFSR
XU19 0 VDD COMP N003 RESET D7 q19 D6 DFFSR
XU20 0 VDD COMP N002 RESET D8 q20 D7 DFFSR
XU21 0 VDD COMP N001 RESET D9 q21 D8 DFFSR
XU23 0 VDD 0 EOC RESET N011 q23 0 DFFSR
.ends SAR

*DAC R-2R

.subckt DAC 1 0 vref D9 D8 D7 D6 D5 D4 D3 D2 D1 D0 out
R1 D9_ out 12k
R2 i out 6k
R3 D8_ i 12k
R4 h i 6k
R5 D7_ h 12k
R6 g h 6k
R7 D6_ g 12k
R8 f g 6k
R9 D5_ f 12k
R10 e f 6k
R11 D4_ e 12k
R12 d e 6k
R13 D3_ d 12k
R14 c d 6k
R15 D2_ c 12k
R16 b c 6k
R17 D1_ b 12k
R18 a b 6k
R19 D0_ a 12k
R20 a 0 12k
X1  D0 D0_ vref 1 0 switch
X2  D1 D1_ vref 1 0 switch
X3  D2 D2_ vref 1 0 switch
X4  D3 D3_ vref 1 0 switch
X5  D4 D4_ vref 1 0 switch
X6  D5 D5_ vref 1 0 switch
X7  D6 D6_ vref 1 0 switch
X8  D7 D7_ vref 1 0 switch
X9  D8 D8_ vref 1 0 switch
X10 D9 D9_ vref 1 0 switch
.ends DAC

.SUBCKT switch data node vref s o
m1t node data_bar vref s pfet W=4u L=0.2u
m2t node data_bar o o nfet W=1u L=0.2u
m3t data_bar data s s pfet W=1.2u L=0.2u
m4t data_bar data o o nfet W=0.6u L=0.2u
.ENDS switch

******************************************

X1 1 0 in clk1 out_sam sample
X2 1 1d 0 out_sam out_dac out_comp comparator
X3 1d 0 clk clk1 clkdivider
X4 1d 0 SOC clk out_comp D9 D8 D7 D6 D5 D4 D3 D2 D1 D0 EOC SAR
X5 1 0 vref D9 D8 D7 D6 D5 D4 D3 D2 D1 D0 out_dac DAC
*************************************

V_a 1 0 3.3v
V_d 1d 0 1.8V
V_ref vref 0 3.3V
V_soc SOC 0 PULSE(0 1.8 1ns 1ns 1ns 0.5us 6us)
V_clk clk 0 PULSE(0 1.8 1n 1n 1n 0.25u 0.5u)
*************************************
*Vin in 0 SINE(1.65v 1.65v 5k)

*********CHANGE INPUT HERE*************

Vin in 0 2000mV
*************************************

.tran 1u 15u
.control
run

plot V(D0) V(D1)+2 V(D2)+4 V(D3)+6 V(D4)+8 V(D5)+10 V(D6)+12 V(D7)+14 V(D8)+16 V(D9)+18 V(EOC)+20 V(SOC)+22 V(clk)+24
*set color0=white
.endc
.end




