magic
tech scmos
timestamp 1598176218
<< nwell >>
rect -70 -199 460 -129
<< ntransistor >>
rect -55 -215 -53 -205
rect -35 -211 -33 -205
rect -2 -215 0 -205
rect 18 -211 20 -205
rect 51 -215 53 -205
rect 71 -211 73 -205
rect 104 -215 106 -205
rect 124 -211 126 -205
rect 157 -215 159 -205
rect 177 -211 179 -205
rect 210 -215 212 -205
rect 230 -211 232 -205
rect 263 -215 265 -205
rect 283 -211 285 -205
rect 316 -215 318 -205
rect 336 -211 338 -205
rect 369 -215 371 -205
rect 389 -211 391 -205
rect 422 -215 424 -205
rect 442 -211 444 -205
<< ptransistor >>
rect -55 -193 -53 -153
rect -35 -165 -33 -153
rect -2 -193 0 -153
rect 18 -165 20 -153
rect 51 -193 53 -153
rect 71 -165 73 -153
rect 104 -193 106 -153
rect 124 -165 126 -153
rect 157 -193 159 -153
rect 177 -165 179 -153
rect 210 -193 212 -153
rect 230 -165 232 -153
rect 263 -193 265 -153
rect 283 -165 285 -153
rect 316 -193 318 -153
rect 336 -165 338 -153
rect 369 -193 371 -153
rect 389 -165 391 -153
rect 422 -193 424 -153
rect 442 -165 444 -153
<< ndiffusion >>
rect -56 -215 -55 -205
rect -53 -215 -52 -205
rect -36 -211 -35 -205
rect -33 -211 -32 -205
rect -3 -215 -2 -205
rect 0 -215 1 -205
rect 17 -211 18 -205
rect 20 -211 21 -205
rect 50 -215 51 -205
rect 53 -215 54 -205
rect 70 -211 71 -205
rect 73 -211 74 -205
rect 103 -215 104 -205
rect 106 -215 107 -205
rect 123 -211 124 -205
rect 126 -211 127 -205
rect 156 -215 157 -205
rect 159 -215 160 -205
rect 176 -211 177 -205
rect 179 -211 180 -205
rect 209 -215 210 -205
rect 212 -215 213 -205
rect 229 -211 230 -205
rect 232 -211 233 -205
rect 262 -215 263 -205
rect 265 -215 266 -205
rect 282 -211 283 -205
rect 285 -211 286 -205
rect 315 -215 316 -205
rect 318 -215 319 -205
rect 335 -211 336 -205
rect 338 -211 339 -205
rect 368 -215 369 -205
rect 371 -215 372 -205
rect 388 -211 389 -205
rect 391 -211 392 -205
rect 421 -215 422 -205
rect 424 -215 425 -205
rect 441 -211 442 -205
rect 444 -211 445 -205
<< pdiffusion >>
rect -56 -159 -55 -153
rect -61 -163 -55 -159
rect -56 -169 -55 -163
rect -61 -175 -55 -169
rect -56 -181 -55 -175
rect -61 -187 -55 -181
rect -56 -193 -55 -187
rect -53 -159 -52 -153
rect -53 -163 -47 -159
rect -53 -169 -52 -163
rect -36 -158 -35 -153
rect -41 -160 -35 -158
rect -36 -165 -35 -160
rect -33 -158 -32 -153
rect -33 -160 -27 -158
rect -33 -165 -32 -160
rect -3 -159 -2 -153
rect -8 -163 -2 -159
rect -53 -175 -47 -169
rect -53 -181 -52 -175
rect -53 -187 -47 -181
rect -53 -193 -52 -187
rect -3 -169 -2 -163
rect -8 -175 -2 -169
rect -3 -181 -2 -175
rect -8 -187 -2 -181
rect -3 -193 -2 -187
rect 0 -159 1 -153
rect 0 -163 6 -159
rect 0 -169 1 -163
rect 17 -158 18 -153
rect 12 -160 18 -158
rect 17 -165 18 -160
rect 20 -158 21 -153
rect 20 -160 26 -158
rect 20 -165 21 -160
rect 50 -159 51 -153
rect 45 -163 51 -159
rect 0 -175 6 -169
rect 0 -181 1 -175
rect 0 -187 6 -181
rect 0 -193 1 -187
rect 50 -169 51 -163
rect 45 -175 51 -169
rect 50 -181 51 -175
rect 45 -187 51 -181
rect 50 -193 51 -187
rect 53 -159 54 -153
rect 53 -163 59 -159
rect 53 -169 54 -163
rect 70 -158 71 -153
rect 65 -160 71 -158
rect 70 -165 71 -160
rect 73 -158 74 -153
rect 73 -160 79 -158
rect 73 -165 74 -160
rect 103 -159 104 -153
rect 98 -163 104 -159
rect 53 -175 59 -169
rect 53 -181 54 -175
rect 53 -187 59 -181
rect 53 -193 54 -187
rect 103 -169 104 -163
rect 98 -175 104 -169
rect 103 -181 104 -175
rect 98 -187 104 -181
rect 103 -193 104 -187
rect 106 -159 107 -153
rect 106 -163 112 -159
rect 106 -169 107 -163
rect 123 -158 124 -153
rect 118 -160 124 -158
rect 123 -165 124 -160
rect 126 -158 127 -153
rect 126 -160 132 -158
rect 126 -165 127 -160
rect 156 -159 157 -153
rect 151 -163 157 -159
rect 106 -175 112 -169
rect 106 -181 107 -175
rect 106 -187 112 -181
rect 106 -193 107 -187
rect 156 -169 157 -163
rect 151 -175 157 -169
rect 156 -181 157 -175
rect 151 -187 157 -181
rect 156 -193 157 -187
rect 159 -159 160 -153
rect 159 -163 165 -159
rect 159 -169 160 -163
rect 176 -158 177 -153
rect 171 -160 177 -158
rect 176 -165 177 -160
rect 179 -158 180 -153
rect 179 -160 185 -158
rect 179 -165 180 -160
rect 209 -159 210 -153
rect 204 -163 210 -159
rect 159 -175 165 -169
rect 159 -181 160 -175
rect 159 -187 165 -181
rect 159 -193 160 -187
rect 209 -169 210 -163
rect 204 -175 210 -169
rect 209 -181 210 -175
rect 204 -187 210 -181
rect 209 -193 210 -187
rect 212 -159 213 -153
rect 212 -163 218 -159
rect 212 -169 213 -163
rect 229 -158 230 -153
rect 224 -160 230 -158
rect 229 -165 230 -160
rect 232 -158 233 -153
rect 232 -160 238 -158
rect 232 -165 233 -160
rect 262 -159 263 -153
rect 257 -163 263 -159
rect 212 -175 218 -169
rect 212 -181 213 -175
rect 212 -187 218 -181
rect 212 -193 213 -187
rect 262 -169 263 -163
rect 257 -175 263 -169
rect 262 -181 263 -175
rect 257 -187 263 -181
rect 262 -193 263 -187
rect 265 -159 266 -153
rect 265 -163 271 -159
rect 265 -169 266 -163
rect 282 -158 283 -153
rect 277 -160 283 -158
rect 282 -165 283 -160
rect 285 -158 286 -153
rect 285 -160 291 -158
rect 285 -165 286 -160
rect 315 -159 316 -153
rect 310 -163 316 -159
rect 265 -175 271 -169
rect 265 -181 266 -175
rect 265 -187 271 -181
rect 265 -193 266 -187
rect 315 -169 316 -163
rect 310 -175 316 -169
rect 315 -181 316 -175
rect 310 -187 316 -181
rect 315 -193 316 -187
rect 318 -159 319 -153
rect 318 -163 324 -159
rect 318 -169 319 -163
rect 335 -158 336 -153
rect 330 -160 336 -158
rect 335 -165 336 -160
rect 338 -158 339 -153
rect 338 -160 344 -158
rect 338 -165 339 -160
rect 368 -159 369 -153
rect 363 -163 369 -159
rect 318 -175 324 -169
rect 318 -181 319 -175
rect 318 -187 324 -181
rect 318 -193 319 -187
rect 368 -169 369 -163
rect 363 -175 369 -169
rect 368 -181 369 -175
rect 363 -187 369 -181
rect 368 -193 369 -187
rect 371 -159 372 -153
rect 371 -163 377 -159
rect 371 -169 372 -163
rect 388 -158 389 -153
rect 383 -160 389 -158
rect 388 -165 389 -160
rect 391 -158 392 -153
rect 391 -160 397 -158
rect 391 -165 392 -160
rect 421 -159 422 -153
rect 416 -163 422 -159
rect 371 -175 377 -169
rect 371 -181 372 -175
rect 371 -187 377 -181
rect 371 -193 372 -187
rect 421 -169 422 -163
rect 416 -175 422 -169
rect 421 -181 422 -175
rect 416 -187 422 -181
rect 421 -193 422 -187
rect 424 -159 425 -153
rect 424 -163 430 -159
rect 424 -169 425 -163
rect 441 -158 442 -153
rect 436 -160 442 -158
rect 441 -165 442 -160
rect 444 -158 445 -153
rect 444 -160 450 -158
rect 444 -165 445 -160
rect 424 -175 430 -169
rect 424 -181 425 -175
rect 424 -187 430 -181
rect 424 -193 425 -187
<< ndcontact >>
rect -61 -215 -56 -205
rect -52 -215 -47 -205
rect -41 -211 -36 -205
rect -32 -211 -27 -205
rect -8 -215 -3 -205
rect 1 -215 6 -205
rect 12 -211 17 -205
rect 21 -211 26 -205
rect 45 -215 50 -205
rect 54 -215 59 -205
rect 65 -211 70 -205
rect 74 -211 79 -205
rect 98 -215 103 -205
rect 107 -215 112 -205
rect 118 -211 123 -205
rect 127 -211 132 -205
rect 151 -215 156 -205
rect 160 -215 165 -205
rect 171 -211 176 -205
rect 180 -211 185 -205
rect 204 -215 209 -205
rect 213 -215 218 -205
rect 224 -211 229 -205
rect 233 -211 238 -205
rect 257 -215 262 -205
rect 266 -215 271 -205
rect 277 -211 282 -205
rect 286 -211 291 -205
rect 310 -215 315 -205
rect 319 -215 324 -205
rect 330 -211 335 -205
rect 339 -211 344 -205
rect 363 -215 368 -205
rect 372 -215 377 -205
rect 383 -211 388 -205
rect 392 -211 397 -205
rect 416 -215 421 -205
rect 425 -215 430 -205
rect 436 -211 441 -205
rect 445 -211 450 -205
<< pdcontact >>
rect -61 -159 -56 -153
rect -61 -169 -56 -163
rect -61 -181 -56 -175
rect -61 -193 -56 -187
rect -52 -159 -47 -153
rect -52 -169 -47 -163
rect -41 -158 -36 -153
rect -41 -165 -36 -160
rect -32 -158 -27 -153
rect -32 -165 -27 -160
rect -8 -159 -3 -153
rect -52 -181 -47 -175
rect -52 -193 -47 -187
rect -8 -169 -3 -163
rect -8 -181 -3 -175
rect -8 -193 -3 -187
rect 1 -159 6 -153
rect 1 -169 6 -163
rect 12 -158 17 -153
rect 12 -165 17 -160
rect 21 -158 26 -153
rect 21 -165 26 -160
rect 45 -159 50 -153
rect 1 -181 6 -175
rect 1 -193 6 -187
rect 45 -169 50 -163
rect 45 -181 50 -175
rect 45 -193 50 -187
rect 54 -159 59 -153
rect 54 -169 59 -163
rect 65 -158 70 -153
rect 65 -165 70 -160
rect 74 -158 79 -153
rect 74 -165 79 -160
rect 98 -159 103 -153
rect 54 -181 59 -175
rect 54 -193 59 -187
rect 98 -169 103 -163
rect 98 -181 103 -175
rect 98 -193 103 -187
rect 107 -159 112 -153
rect 107 -169 112 -163
rect 118 -158 123 -153
rect 118 -165 123 -160
rect 127 -158 132 -153
rect 127 -165 132 -160
rect 151 -159 156 -153
rect 107 -181 112 -175
rect 107 -193 112 -187
rect 151 -169 156 -163
rect 151 -181 156 -175
rect 151 -193 156 -187
rect 160 -159 165 -153
rect 160 -169 165 -163
rect 171 -158 176 -153
rect 171 -165 176 -160
rect 180 -158 185 -153
rect 180 -165 185 -160
rect 204 -159 209 -153
rect 160 -181 165 -175
rect 160 -193 165 -187
rect 204 -169 209 -163
rect 204 -181 209 -175
rect 204 -193 209 -187
rect 213 -159 218 -153
rect 213 -169 218 -163
rect 224 -158 229 -153
rect 224 -165 229 -160
rect 233 -158 238 -153
rect 233 -165 238 -160
rect 257 -159 262 -153
rect 213 -181 218 -175
rect 213 -193 218 -187
rect 257 -169 262 -163
rect 257 -181 262 -175
rect 257 -193 262 -187
rect 266 -159 271 -153
rect 266 -169 271 -163
rect 277 -158 282 -153
rect 277 -165 282 -160
rect 286 -158 291 -153
rect 286 -165 291 -160
rect 310 -159 315 -153
rect 266 -181 271 -175
rect 266 -193 271 -187
rect 310 -169 315 -163
rect 310 -181 315 -175
rect 310 -193 315 -187
rect 319 -159 324 -153
rect 319 -169 324 -163
rect 330 -158 335 -153
rect 330 -165 335 -160
rect 339 -158 344 -153
rect 339 -165 344 -160
rect 363 -159 368 -153
rect 319 -181 324 -175
rect 319 -193 324 -187
rect 363 -169 368 -163
rect 363 -181 368 -175
rect 363 -193 368 -187
rect 372 -159 377 -153
rect 372 -169 377 -163
rect 383 -158 388 -153
rect 383 -165 388 -160
rect 392 -158 397 -153
rect 392 -165 397 -160
rect 416 -159 421 -153
rect 372 -181 377 -175
rect 372 -193 377 -187
rect 416 -169 421 -163
rect 416 -181 421 -175
rect 416 -193 421 -187
rect 425 -159 430 -153
rect 425 -169 430 -163
rect 436 -158 441 -153
rect 436 -165 441 -160
rect 445 -158 450 -153
rect 445 -165 450 -160
rect 425 -181 430 -175
rect 425 -193 430 -187
<< psubstratepcontact >>
rect -67 -229 -63 -223
rect -56 -229 -52 -223
rect -44 -229 -40 -223
rect -34 -229 -30 -223
rect -25 -229 -21 -223
rect -14 -229 -10 -223
rect -3 -229 1 -223
rect 9 -229 13 -223
rect 19 -229 23 -223
rect 28 -229 32 -223
rect 39 -229 43 -223
rect 50 -229 54 -223
rect 62 -229 66 -223
rect 72 -229 76 -223
rect 81 -229 85 -223
rect 92 -229 96 -223
rect 103 -229 107 -223
rect 115 -229 119 -223
rect 125 -229 129 -223
rect 134 -229 138 -223
rect 145 -229 149 -223
rect 156 -229 160 -223
rect 168 -229 172 -223
rect 178 -229 182 -223
rect 187 -229 191 -223
rect 198 -229 202 -223
rect 209 -229 213 -223
rect 221 -229 225 -223
rect 231 -229 235 -223
rect 240 -229 244 -223
rect 251 -229 255 -223
rect 262 -229 266 -223
rect 274 -229 278 -223
rect 284 -229 288 -223
rect 293 -229 297 -223
rect 304 -229 308 -223
rect 315 -229 319 -223
rect 327 -229 331 -223
rect 337 -229 341 -223
rect 346 -229 350 -223
rect 357 -229 361 -223
rect 368 -229 372 -223
rect 380 -229 384 -223
rect 390 -229 394 -223
rect 399 -229 403 -223
rect 410 -229 414 -223
rect 421 -229 425 -223
rect 433 -229 437 -223
rect 443 -229 447 -223
rect 452 -229 456 -223
<< nsubstratencontact >>
rect 1 85 13 91
rect 1 1 13 7
rect 21 85 33 91
rect 21 1 33 7
rect 41 85 53 91
rect 41 1 53 7
rect 81 85 93 91
rect 81 1 93 7
rect 101 85 113 91
rect 101 1 113 7
rect 121 85 133 91
rect 121 1 133 7
rect 161 85 173 91
rect 161 1 173 7
rect 181 85 193 91
rect 181 1 193 7
rect 201 85 213 91
rect 201 1 213 7
rect 241 85 253 91
rect 241 1 253 7
rect 261 85 273 91
rect 261 1 273 7
rect 281 85 293 91
rect 281 1 293 7
rect 321 85 333 91
rect 321 1 333 7
rect 341 85 353 91
rect 341 1 353 7
rect 361 85 373 91
rect 361 1 373 7
rect 1 -16 13 -10
rect 1 -100 13 -94
rect 41 -15 53 -9
rect 41 -99 53 -93
rect 61 -15 73 -9
rect 61 -99 73 -93
rect 81 -15 93 -9
rect 81 -99 93 -93
rect 121 -15 133 -9
rect 121 -99 133 -93
rect 141 -15 153 -9
rect 141 -99 153 -93
rect 161 -15 173 -9
rect 161 -99 173 -93
rect 201 -15 213 -9
rect 201 -99 213 -93
rect 221 -15 233 -9
rect 221 -99 233 -93
rect 241 -15 253 -9
rect 241 -99 253 -93
rect 281 -15 293 -9
rect 281 -99 293 -93
rect 301 -15 313 -9
rect 301 -99 313 -93
rect 321 -15 333 -9
rect 321 -99 333 -93
rect 361 -15 373 -9
rect 361 -99 373 -93
rect 381 -15 393 -9
rect 381 -99 393 -93
rect -67 -139 -63 -133
rect -57 -139 -53 -133
rect -48 -139 -44 -133
rect -40 -139 -36 -133
rect -32 -139 -28 -133
rect -24 -139 -20 -133
rect -14 -139 -10 -133
rect -4 -139 0 -133
rect 5 -139 9 -133
rect 13 -139 17 -133
rect 21 -139 25 -133
rect 29 -139 33 -133
rect 39 -139 43 -133
rect 49 -139 53 -133
rect 58 -139 62 -133
rect 66 -139 70 -133
rect 74 -139 78 -133
rect 82 -139 86 -133
rect 92 -139 96 -133
rect 102 -139 106 -133
rect 111 -139 115 -133
rect 119 -139 123 -133
rect 127 -139 131 -133
rect 135 -139 139 -133
rect 145 -139 149 -133
rect 155 -139 159 -133
rect 164 -139 168 -133
rect 172 -139 176 -133
rect 180 -139 184 -133
rect 188 -139 192 -133
rect 198 -139 202 -133
rect 208 -139 212 -133
rect 217 -139 221 -133
rect 225 -139 229 -133
rect 233 -139 237 -133
rect 241 -139 245 -133
rect 251 -139 255 -133
rect 261 -139 265 -133
rect 270 -139 274 -133
rect 278 -139 282 -133
rect 286 -139 290 -133
rect 294 -139 298 -133
rect 304 -139 308 -133
rect 314 -139 318 -133
rect 323 -139 327 -133
rect 331 -139 335 -133
rect 339 -139 343 -133
rect 347 -139 351 -133
rect 357 -139 361 -133
rect 367 -139 371 -133
rect 376 -139 380 -133
rect 384 -139 388 -133
rect 392 -139 396 -133
rect 400 -139 404 -133
rect 410 -139 414 -133
rect 420 -139 424 -133
rect 429 -139 433 -133
rect 437 -139 441 -133
rect 445 -139 449 -133
rect 453 -139 457 -133
<< polysilicon >>
rect -55 -147 -31 -143
rect -2 -147 22 -143
rect 51 -147 75 -143
rect 104 -147 128 -143
rect 157 -147 181 -143
rect 210 -147 234 -143
rect 263 -147 287 -143
rect 316 -147 340 -143
rect 369 -147 393 -143
rect 422 -147 446 -143
rect -55 -153 -53 -147
rect -35 -153 -33 -150
rect -2 -153 0 -147
rect 18 -153 20 -150
rect 51 -153 53 -147
rect 71 -153 73 -150
rect 104 -153 106 -147
rect 124 -153 126 -150
rect 157 -153 159 -147
rect 177 -153 179 -150
rect 210 -153 212 -147
rect 230 -153 232 -150
rect 263 -153 265 -147
rect 283 -153 285 -150
rect 316 -153 318 -147
rect 336 -153 338 -150
rect 369 -153 371 -147
rect 389 -153 391 -150
rect 422 -153 424 -147
rect 442 -153 444 -150
rect -55 -205 -53 -193
rect -35 -205 -33 -165
rect -2 -205 0 -193
rect 18 -205 20 -165
rect 51 -205 53 -193
rect 71 -205 73 -165
rect 104 -205 106 -193
rect 124 -205 126 -165
rect 157 -205 159 -193
rect 177 -205 179 -165
rect 210 -205 212 -193
rect 230 -205 232 -165
rect 263 -205 265 -193
rect 283 -205 285 -165
rect 316 -205 318 -193
rect 336 -205 338 -165
rect 369 -205 371 -193
rect 389 -205 391 -165
rect 422 -205 424 -193
rect 442 -205 444 -165
rect -35 -214 -33 -211
rect -55 -218 -53 -215
rect -2 -218 0 -215
rect 18 -218 20 -211
rect 51 -218 53 -215
rect 71 -218 73 -211
rect 104 -218 106 -215
rect 124 -218 126 -211
rect 157 -218 159 -215
rect 177 -218 179 -211
rect 210 -218 212 -215
rect 230 -218 232 -211
rect 263 -218 265 -215
rect 283 -218 285 -211
rect 316 -218 318 -215
rect 336 -218 338 -211
rect 369 -218 371 -215
rect 389 -218 391 -211
rect 422 -218 424 -215
rect 442 -218 444 -211
<< polycontact >>
rect -31 -147 -27 -143
rect 22 -147 26 -143
rect 75 -147 79 -143
rect 128 -147 132 -143
rect 181 -147 185 -143
rect 234 -147 238 -143
rect 287 -147 291 -143
rect 340 -147 344 -143
rect 393 -147 397 -143
rect 446 -147 450 -143
<< metal1 >>
rect 45 91 49 94
rect 125 91 129 94
rect 205 91 209 94
rect 285 91 289 94
rect 365 91 369 94
rect -12 85 1 91
rect 13 85 21 91
rect 65 85 81 91
rect 93 85 101 91
rect 145 85 161 91
rect 173 85 181 91
rect 225 85 241 91
rect 253 85 261 91
rect 305 85 321 91
rect 333 85 341 91
rect 5 -10 9 1
rect 25 -93 29 1
rect 45 -9 49 1
rect 65 -9 69 85
rect 85 -9 89 1
rect 105 -93 109 1
rect 125 -9 129 1
rect 145 -9 149 85
rect 165 -9 169 1
rect 185 -93 189 1
rect 205 -9 209 1
rect 225 -9 229 85
rect 245 -9 249 1
rect 265 -93 269 1
rect 285 -9 289 1
rect 305 -9 309 85
rect 325 -9 329 1
rect 345 -93 349 1
rect 365 -9 369 1
rect 385 -9 389 -4
rect 25 -99 41 -93
rect 53 -99 61 -93
rect 105 -99 121 -93
rect 133 -99 141 -93
rect 185 -99 201 -93
rect 213 -99 221 -93
rect 265 -99 281 -93
rect 293 -99 301 -93
rect 345 -99 361 -93
rect 373 -99 381 -93
rect 5 -107 9 -100
rect 85 -106 89 -99
rect 165 -110 169 -99
rect 245 -106 249 -99
rect 325 -106 329 -99
rect -70 -133 460 -132
rect -70 -139 -67 -133
rect -63 -139 -57 -133
rect -53 -139 -48 -133
rect -44 -139 -40 -133
rect -36 -139 -32 -133
rect -28 -139 -24 -133
rect -20 -139 -14 -133
rect -10 -139 -4 -133
rect 0 -139 5 -133
rect 9 -139 13 -133
rect 17 -139 21 -133
rect 25 -139 29 -133
rect 33 -139 39 -133
rect 43 -139 49 -133
rect 53 -139 58 -133
rect 62 -139 66 -133
rect 70 -139 74 -133
rect 78 -139 82 -133
rect 86 -139 92 -133
rect 96 -139 102 -133
rect 106 -139 111 -133
rect 115 -139 119 -133
rect 123 -139 127 -133
rect 131 -139 135 -133
rect 139 -139 145 -133
rect 149 -139 155 -133
rect 159 -139 164 -133
rect 168 -139 172 -133
rect 176 -139 180 -133
rect 184 -139 188 -133
rect 192 -139 198 -133
rect 202 -139 208 -133
rect 212 -139 217 -133
rect 221 -139 225 -133
rect 229 -139 233 -133
rect 237 -139 241 -133
rect 245 -139 251 -133
rect 255 -139 261 -133
rect 265 -139 270 -133
rect 274 -139 278 -133
rect 282 -139 286 -133
rect 290 -139 294 -133
rect 298 -139 304 -133
rect 308 -139 314 -133
rect 318 -139 323 -133
rect 327 -139 331 -133
rect 335 -139 339 -133
rect 343 -139 347 -133
rect 351 -139 357 -133
rect 361 -139 367 -133
rect 371 -139 376 -133
rect 380 -139 384 -133
rect 388 -139 392 -133
rect 396 -139 400 -133
rect 404 -139 410 -133
rect 414 -139 420 -133
rect 424 -139 429 -133
rect 433 -139 437 -133
rect 441 -139 445 -133
rect 449 -139 453 -133
rect 457 -139 460 -133
rect -70 -140 460 -139
rect -41 -153 -36 -140
rect -31 -153 -27 -147
rect 12 -153 17 -140
rect 22 -153 26 -147
rect 65 -153 70 -140
rect 75 -153 79 -147
rect 118 -153 123 -140
rect 128 -153 132 -147
rect 171 -153 176 -140
rect 181 -153 185 -147
rect 224 -153 229 -140
rect 234 -153 238 -147
rect 277 -153 282 -140
rect 287 -153 291 -147
rect 330 -153 335 -140
rect 340 -153 344 -147
rect 383 -153 388 -140
rect 393 -153 397 -147
rect 436 -153 441 -140
rect 446 -153 450 -147
rect -61 -163 -56 -159
rect -61 -175 -56 -169
rect -61 -187 -56 -181
rect -82 -199 -76 -193
rect -52 -163 -47 -159
rect -41 -160 -36 -158
rect -32 -160 -27 -158
rect -52 -175 -47 -169
rect -52 -187 -47 -181
rect -52 -205 -47 -193
rect -32 -205 -27 -165
rect -8 -163 -3 -159
rect -8 -175 -3 -169
rect -8 -187 -3 -181
rect 1 -163 6 -159
rect 12 -160 17 -158
rect 21 -160 26 -158
rect 1 -175 6 -169
rect 1 -187 6 -181
rect 1 -205 6 -193
rect 21 -205 26 -165
rect 45 -163 50 -159
rect 45 -175 50 -169
rect 45 -187 50 -181
rect 54 -163 59 -159
rect 65 -160 70 -158
rect 74 -160 79 -158
rect 54 -175 59 -169
rect 54 -187 59 -181
rect 54 -205 59 -193
rect 74 -205 79 -165
rect 98 -163 103 -159
rect 98 -175 103 -169
rect 98 -187 103 -181
rect 107 -163 112 -159
rect 118 -160 123 -158
rect 127 -160 132 -158
rect 107 -175 112 -169
rect 107 -187 112 -181
rect 107 -205 112 -193
rect 127 -205 132 -165
rect 151 -163 156 -159
rect 151 -175 156 -169
rect 151 -187 156 -181
rect 160 -163 165 -159
rect 171 -160 176 -158
rect 180 -160 185 -158
rect 160 -175 165 -169
rect 160 -187 165 -181
rect 160 -205 165 -193
rect 180 -205 185 -165
rect 204 -163 209 -159
rect 204 -175 209 -169
rect 204 -187 209 -181
rect 213 -163 218 -159
rect 224 -160 229 -158
rect 233 -160 238 -158
rect 213 -175 218 -169
rect 213 -187 218 -181
rect 213 -205 218 -193
rect 233 -205 238 -165
rect 257 -163 262 -159
rect 257 -175 262 -169
rect 257 -187 262 -181
rect 266 -163 271 -159
rect 277 -160 282 -158
rect 286 -160 291 -158
rect 266 -175 271 -169
rect 266 -187 271 -181
rect 266 -205 271 -193
rect 286 -205 291 -165
rect 310 -163 315 -159
rect 310 -175 315 -169
rect 310 -187 315 -181
rect 319 -163 324 -159
rect 330 -160 335 -158
rect 339 -160 344 -158
rect 319 -175 324 -169
rect 319 -187 324 -181
rect 319 -205 324 -193
rect 339 -205 344 -165
rect 363 -163 368 -159
rect 363 -175 368 -169
rect 363 -187 368 -181
rect 372 -163 377 -159
rect 383 -160 388 -158
rect 392 -160 397 -158
rect 372 -175 377 -169
rect 372 -187 377 -181
rect 372 -205 377 -193
rect 392 -205 397 -165
rect 416 -163 421 -159
rect 416 -175 421 -169
rect 416 -187 421 -181
rect 425 -163 430 -159
rect 436 -160 441 -158
rect 445 -160 450 -158
rect 425 -175 430 -169
rect 425 -187 430 -181
rect 425 -205 430 -193
rect 445 -205 450 -165
rect -61 -222 -56 -215
rect -41 -222 -36 -211
rect -8 -222 -3 -215
rect 12 -222 17 -211
rect 45 -222 50 -215
rect 65 -222 70 -211
rect 98 -222 103 -215
rect 118 -222 123 -211
rect 151 -222 156 -215
rect 171 -222 176 -211
rect 204 -222 209 -215
rect 224 -222 229 -211
rect 257 -222 262 -215
rect 277 -222 282 -211
rect 310 -222 315 -215
rect 330 -222 335 -211
rect 363 -222 368 -215
rect 383 -222 388 -211
rect 416 -222 421 -215
rect 436 -222 441 -211
rect 460 -222 465 -205
rect -70 -223 465 -222
rect -70 -229 -67 -223
rect -63 -229 -56 -223
rect -52 -229 -44 -223
rect -40 -229 -34 -223
rect -30 -229 -25 -223
rect -21 -229 -14 -223
rect -10 -229 -3 -223
rect 1 -229 9 -223
rect 13 -229 19 -223
rect 23 -229 28 -223
rect 32 -229 39 -223
rect 43 -229 50 -223
rect 54 -229 62 -223
rect 66 -229 72 -223
rect 76 -229 81 -223
rect 85 -229 92 -223
rect 96 -229 103 -223
rect 107 -229 115 -223
rect 119 -229 125 -223
rect 129 -229 134 -223
rect 138 -229 145 -223
rect 149 -229 156 -223
rect 160 -229 168 -223
rect 172 -229 178 -223
rect 182 -229 187 -223
rect 191 -229 198 -223
rect 202 -229 209 -223
rect 213 -229 221 -223
rect 225 -229 231 -223
rect 235 -229 240 -223
rect 244 -229 251 -223
rect 255 -229 262 -223
rect 266 -229 274 -223
rect 278 -229 284 -223
rect 288 -229 293 -223
rect 297 -229 304 -223
rect 308 -229 315 -223
rect 319 -229 327 -223
rect 331 -229 337 -223
rect 341 -229 346 -223
rect 350 -229 357 -223
rect 361 -229 368 -223
rect 372 -229 380 -223
rect 384 -229 390 -223
rect 394 -229 399 -223
rect 403 -229 410 -223
rect 414 -229 421 -223
rect 425 -229 433 -223
rect 437 -229 443 -223
rect 447 -229 452 -223
rect 456 -229 465 -223
rect -70 -230 465 -229
<< m2contact >>
rect 45 94 49 98
rect 125 94 129 98
rect 205 94 209 98
rect 285 94 289 98
rect 365 94 369 98
rect 385 -4 389 1
rect 5 -111 9 -107
rect 85 -110 89 -106
rect 160 -110 165 -106
rect 245 -110 249 -106
rect 325 -110 329 -106
rect -76 -199 -71 -193
rect -61 -199 -56 -193
rect -52 -159 -47 -153
rect -8 -199 -3 -193
rect 1 -159 6 -153
rect 45 -199 50 -193
rect 54 -159 59 -153
rect 98 -199 103 -193
rect 107 -159 112 -153
rect 151 -199 156 -193
rect 160 -159 165 -153
rect 204 -199 209 -193
rect 213 -159 218 -153
rect 257 -199 262 -193
rect 266 -159 271 -153
rect 310 -199 315 -193
rect 319 -159 324 -153
rect 363 -199 368 -193
rect 372 -159 377 -153
rect 416 -199 421 -193
rect 425 -159 430 -153
rect 460 -205 465 -199
<< metal2 >>
rect -52 -111 5 -107
rect -52 -153 -47 -111
rect 45 -116 49 94
rect 1 -121 49 -116
rect 54 -110 85 -106
rect 125 -110 129 94
rect 205 -106 209 94
rect 1 -153 6 -121
rect 54 -153 59 -110
rect 107 -115 129 -110
rect 205 -110 218 -106
rect 249 -110 271 -106
rect 107 -153 112 -115
rect 160 -153 165 -110
rect 213 -153 218 -110
rect 266 -153 271 -110
rect 285 -116 289 94
rect 365 -105 369 94
rect 389 -4 465 1
rect 329 -110 343 -106
rect 365 -109 430 -105
rect 285 -121 324 -116
rect 319 -153 324 -121
rect 339 -120 343 -110
rect 339 -124 377 -120
rect 372 -153 377 -124
rect 425 -153 430 -109
rect -71 -199 -61 -193
rect -56 -199 -8 -193
rect -3 -199 45 -193
rect 50 -199 98 -193
rect 103 -199 151 -193
rect 156 -199 204 -193
rect 209 -199 257 -193
rect 262 -199 310 -193
rect 315 -199 363 -193
rect 368 -199 416 -193
rect 421 -199 449 -193
rect 460 -199 465 -4
<< pseudo_rnwell >>
rect 0 91 14 92
rect 0 1 1 91
rect 13 1 14 91
rect 0 0 14 1
rect 20 91 34 92
rect 20 1 21 91
rect 33 1 34 91
rect 20 0 34 1
rect 40 91 54 92
rect 40 1 41 91
rect 53 1 54 91
rect 40 0 54 1
rect 80 91 94 92
rect 80 1 81 91
rect 93 1 94 91
rect 80 0 94 1
rect 100 91 114 92
rect 100 1 101 91
rect 113 1 114 91
rect 100 0 114 1
rect 120 91 134 92
rect 120 1 121 91
rect 133 1 134 91
rect 120 0 134 1
rect 160 91 174 92
rect 160 1 161 91
rect 173 1 174 91
rect 160 0 174 1
rect 180 91 194 92
rect 180 1 181 91
rect 193 1 194 91
rect 180 0 194 1
rect 200 91 214 92
rect 200 1 201 91
rect 213 1 214 91
rect 200 0 214 1
rect 240 91 254 92
rect 240 1 241 91
rect 253 1 254 91
rect 240 0 254 1
rect 260 91 274 92
rect 260 1 261 91
rect 273 1 274 91
rect 260 0 274 1
rect 280 91 294 92
rect 280 1 281 91
rect 293 1 294 91
rect 280 0 294 1
rect 320 91 334 92
rect 320 1 321 91
rect 333 1 334 91
rect 320 0 334 1
rect 340 91 354 92
rect 340 1 341 91
rect 353 1 354 91
rect 340 0 354 1
rect 360 91 374 92
rect 360 1 361 91
rect 373 1 374 91
rect 360 0 374 1
rect 40 -9 54 -8
rect 0 -10 14 -9
rect 0 -100 1 -10
rect 13 -100 14 -10
rect 40 -99 41 -9
rect 53 -99 54 -9
rect 40 -100 54 -99
rect 60 -9 74 -8
rect 60 -99 61 -9
rect 73 -99 74 -9
rect 60 -100 74 -99
rect 80 -9 94 -8
rect 80 -99 81 -9
rect 93 -99 94 -9
rect 80 -100 94 -99
rect 120 -9 134 -8
rect 120 -99 121 -9
rect 133 -99 134 -9
rect 120 -100 134 -99
rect 140 -9 154 -8
rect 140 -99 141 -9
rect 153 -99 154 -9
rect 140 -100 154 -99
rect 160 -9 174 -8
rect 160 -99 161 -9
rect 173 -99 174 -9
rect 160 -100 174 -99
rect 200 -9 214 -8
rect 200 -99 201 -9
rect 213 -99 214 -9
rect 200 -100 214 -99
rect 220 -9 234 -8
rect 220 -99 221 -9
rect 233 -99 234 -9
rect 220 -100 234 -99
rect 240 -9 254 -8
rect 240 -99 241 -9
rect 253 -99 254 -9
rect 240 -100 254 -99
rect 280 -9 294 -8
rect 280 -99 281 -9
rect 293 -99 294 -9
rect 280 -100 294 -99
rect 300 -9 314 -8
rect 300 -99 301 -9
rect 313 -99 314 -9
rect 300 -100 314 -99
rect 320 -9 334 -8
rect 320 -99 321 -9
rect 333 -99 334 -9
rect 320 -100 334 -99
rect 360 -9 374 -8
rect 360 -99 361 -9
rect 373 -99 374 -9
rect 360 -100 374 -99
rect 380 -9 394 -8
rect 380 -99 381 -9
rect 393 -99 394 -9
rect 380 -100 394 -99
rect 0 -101 14 -100
<< rnwell >>
rect 1 7 13 85
rect 21 7 33 85
rect 41 7 53 85
rect 81 7 93 85
rect 101 7 113 85
rect 121 7 133 85
rect 161 7 173 85
rect 181 7 193 85
rect 201 7 213 85
rect 241 7 253 85
rect 261 7 273 85
rect 281 7 293 85
rect 321 7 333 85
rect 341 7 353 85
rect 361 7 373 85
rect 1 -94 13 -16
rect 41 -93 53 -15
rect 61 -93 73 -15
rect 81 -93 93 -15
rect 121 -93 133 -15
rect 141 -93 153 -15
rect 161 -93 173 -15
rect 201 -93 213 -15
rect 221 -93 233 -15
rect 241 -93 253 -15
rect 281 -93 293 -15
rect 301 -93 313 -15
rect 321 -93 333 -15
rect 361 -93 373 -15
rect 381 -93 393 -15
<< labels >>
rlabel polysilicon -34 -151 -34 -151 1 d9
rlabel polysilicon 19 -152 19 -152 1 d8
rlabel polysilicon 72 -152 72 -152 1 d7
rlabel polysilicon 125 -151 125 -151 1 d6
rlabel polysilicon 178 -151 178 -151 1 d5
rlabel polysilicon 231 -152 231 -152 1 d4
rlabel polysilicon 284 -151 284 -151 1 d3
rlabel polysilicon 337 -152 337 -152 1 d2
rlabel polysilicon 390 -151 390 -151 1 d1
rlabel polysilicon 443 -151 443 -151 1 d0
rlabel metal1 -59 -136 -59 -136 1 1
rlabel metal1 -48 -226 -48 -226 1 0
rlabel metal1 -10 88 -10 88 1 out_dac
rlabel metal1 -79 -196 -79 -196 3 vref
<< end >>
