magic
tech scmos
timestamp 1598189956
<< nwell >>
rect 222 106 229 108
rect 451 106 457 108
rect 679 106 685 108
rect 907 106 916 108
rect 216 100 233 106
rect 445 100 461 106
rect 673 100 689 106
rect 901 100 920 106
rect 222 71 229 100
rect 451 71 457 100
rect 679 71 685 100
rect 907 71 916 100
rect -2 -21 4 -19
rect 226 -21 232 -19
rect 454 -21 460 -19
rect 682 -21 688 -19
rect 910 -21 916 -19
rect -6 -27 10 -21
rect 222 -27 238 -21
rect 450 -27 466 -21
rect 678 -27 694 -21
rect 906 -27 922 -21
rect -2 -56 4 -27
rect 226 -56 232 -27
rect 454 -56 460 -27
rect 682 -53 688 -27
rect 910 -56 916 -27
rect -2 -147 4 -145
rect 226 -147 232 -145
rect 454 -147 460 -145
rect 682 -147 688 -145
rect -8 -153 8 -147
rect 220 -153 236 -147
rect 448 -153 464 -147
rect 676 -153 692 -147
rect -2 -182 4 -153
rect 226 -158 232 -153
rect 226 -174 234 -158
rect 226 -182 232 -174
rect 454 -182 460 -153
rect 682 -182 688 -153
rect 910 -182 916 -145
rect 919 -158 923 -155
rect 919 -166 923 -162
rect 919 -182 923 -171
rect 226 -302 232 -265
rect 454 -302 460 -265
rect 682 -267 688 -265
rect 910 -267 916 -265
rect 678 -273 694 -267
rect 906 -273 922 -267
rect 678 -290 681 -282
rect 682 -290 688 -273
rect 678 -294 688 -290
rect 682 -302 688 -294
rect 905 -295 909 -291
rect 910 -302 916 -273
<< metal1 >>
rect 216 100 233 106
rect 445 100 461 106
rect 673 100 689 106
rect 901 100 920 106
rect 1132 100 1157 106
rect 2 63 3 67
rect 445 63 460 67
rect 673 63 688 67
rect 902 63 919 67
rect 217 54 225 58
rect 446 54 453 58
rect 674 54 681 58
rect 902 54 909 58
rect 1133 54 1168 58
rect -19 50 3 54
rect -19 6 -15 50
rect 221 44 225 54
rect 449 44 453 54
rect 677 44 681 54
rect 905 44 909 54
rect 916 50 919 54
rect -10 40 3 44
rect 221 40 232 44
rect 453 40 460 44
rect 681 40 688 44
rect 909 40 919 44
rect -10 6 -6 40
rect 210 6 214 26
rect 441 6 445 9
rect 669 6 674 9
rect 897 7 898 11
rect 897 6 902 7
rect -19 0 3 6
rect 216 0 232 6
rect 445 0 460 6
rect 673 0 688 6
rect 901 0 919 6
rect -6 -27 10 -21
rect 222 -27 238 -21
rect 450 -27 466 -21
rect 678 -27 694 -21
rect 906 -27 922 -21
rect 1134 -27 1157 -21
rect -231 -73 -219 -69
rect 2 -73 9 -69
rect 230 -73 237 -69
rect 458 -73 465 -69
rect 686 -73 693 -69
rect -230 -186 -226 -73
rect 2 -83 6 -73
rect 230 -83 234 -73
rect 458 -83 462 -73
rect 686 -83 690 -73
rect 914 -83 918 -69
rect 1164 -83 1168 54
rect -5 -87 2 -83
rect 223 -87 234 -83
rect 451 -87 462 -83
rect 679 -87 690 -83
rect 907 -87 918 -83
rect 1135 -87 1164 -83
rect 230 -94 234 -87
rect 458 -95 462 -87
rect -13 -121 -9 -102
rect 215 -121 219 -102
rect 686 -95 690 -87
rect 905 -94 914 -90
rect 443 -121 447 -102
rect 671 -121 675 -103
rect 899 -121 903 -103
rect 1127 -108 1131 -103
rect 1130 -121 1131 -108
rect -5 -127 10 -121
rect 223 -127 238 -121
rect 451 -127 466 -121
rect 679 -127 694 -121
rect 907 -127 922 -121
rect 1135 -127 1149 -121
rect -8 -153 8 -147
rect 220 -153 236 -147
rect 448 -153 464 -147
rect 676 -153 692 -147
rect 904 -153 920 -147
rect 1132 -153 1157 -147
rect 918 -186 922 -183
rect -230 -190 -221 -186
rect 6 -190 7 -186
rect 234 -190 237 -186
rect 462 -190 463 -186
rect 690 -190 691 -186
rect 918 -190 919 -186
rect -7 -199 0 -195
rect 221 -199 228 -195
rect 449 -199 456 -195
rect 677 -199 684 -195
rect 905 -199 912 -195
rect 1132 -199 1152 -195
rect -220 -253 -216 -199
rect -4 -216 0 -199
rect 8 -203 10 -199
rect -4 -220 7 -216
rect 224 -220 228 -199
rect 232 -220 235 -216
rect 452 -220 456 -199
rect 460 -220 463 -216
rect 680 -220 684 -199
rect 694 -213 696 -209
rect 688 -220 691 -216
rect 908 -220 912 -199
rect 916 -220 919 -216
rect -8 -253 7 -247
rect 219 -253 235 -247
rect 447 -253 463 -247
rect 676 -253 691 -247
rect 903 -253 919 -247
rect 222 -273 238 -267
rect 450 -273 466 -267
rect 678 -273 694 -267
rect 906 -273 922 -267
rect 221 -310 225 -302
rect 449 -310 453 -303
rect 677 -310 681 -303
rect 905 -310 909 -303
rect 1138 -310 1145 -306
rect 1 -319 9 -315
rect 230 -319 237 -315
rect 458 -319 465 -315
rect 686 -319 693 -315
rect 914 -319 920 -315
rect 1 -391 5 -319
rect 230 -336 234 -319
rect 458 -336 462 -319
rect 686 -336 690 -319
rect 914 -336 918 -319
rect 1135 -333 1140 -329
rect 1148 -336 1152 -199
rect 223 -340 237 -336
rect 451 -340 462 -336
rect 679 -340 690 -336
rect 907 -340 918 -336
rect 1135 -340 1167 -336
rect 1133 -367 1137 -361
rect 223 -373 238 -367
rect 451 -373 466 -367
rect 679 -373 694 -367
rect 907 -373 922 -367
rect 1135 -373 1155 -367
rect 1163 -392 1167 -340
<< m2contact >>
rect 1157 100 1161 106
rect -2 63 2 67
rect 228 63 232 67
rect 441 63 445 67
rect 669 63 673 67
rect 898 63 902 67
rect 236 50 240 54
rect 463 50 467 54
rect 685 50 689 54
rect 912 50 916 54
rect 449 40 453 44
rect 677 40 681 44
rect 905 40 909 44
rect -1 33 3 37
rect 221 36 225 40
rect 231 33 235 37
rect 456 33 460 37
rect 685 33 689 37
rect 918 33 922 37
rect 210 26 214 30
rect 441 9 445 13
rect 669 9 673 13
rect 898 7 902 11
rect 1132 0 1137 6
rect 1157 -27 1161 -21
rect -5 -77 -1 -73
rect 223 -77 227 -73
rect 451 -77 455 -73
rect 678 -77 682 -73
rect 907 -77 911 -73
rect 918 -73 922 -69
rect 1135 -78 1139 -73
rect 2 -87 6 -83
rect 1164 -87 1168 -83
rect -5 -94 -1 -90
rect 223 -94 227 -90
rect 451 -94 455 -90
rect 230 -98 234 -94
rect 678 -94 682 -90
rect -13 -102 -9 -98
rect 215 -102 219 -98
rect 443 -102 447 -98
rect 458 -99 462 -95
rect 914 -94 918 -90
rect 1135 -94 1139 -90
rect 686 -99 690 -95
rect 671 -103 675 -99
rect 899 -103 903 -99
rect 1127 -103 1131 -99
rect 1149 -127 1153 -121
rect 1157 -153 1161 -147
rect 918 -183 922 -179
rect 2 -190 6 -186
rect 230 -190 234 -186
rect 458 -190 462 -186
rect 686 -190 690 -186
rect 4 -203 8 -199
rect 6 -213 10 -209
rect 233 -203 237 -199
rect 234 -213 238 -209
rect 228 -220 232 -216
rect 461 -203 465 -199
rect 462 -213 466 -209
rect 456 -220 460 -216
rect 688 -203 692 -199
rect 690 -213 694 -209
rect 684 -220 688 -216
rect 916 -203 920 -199
rect 918 -213 922 -209
rect 912 -220 916 -216
rect 1132 -253 1137 -247
rect 1134 -273 1138 -267
rect 221 -302 225 -298
rect 449 -303 453 -299
rect 677 -303 681 -299
rect 905 -303 909 -299
rect 1134 -310 1138 -306
rect 466 -319 470 -315
rect 693 -319 697 -315
rect 920 -319 924 -315
rect 222 -323 226 -319
rect 221 -333 225 -329
rect 451 -323 455 -319
rect 448 -333 452 -329
rect 676 -323 680 -319
rect 676 -333 680 -329
rect 906 -323 910 -319
rect 905 -333 909 -329
rect 1133 -323 1137 -319
rect 1140 -333 1144 -329
rect 237 -340 241 -336
rect 1133 -361 1137 -357
rect 1155 -373 1159 -367
<< metal2 >>
rect -10 63 -2 67
rect 2 63 7 67
rect 210 63 228 67
rect -1 -3 3 33
rect 210 30 214 63
rect 233 50 236 54
rect 221 31 225 36
rect 231 -3 235 33
rect 441 13 445 63
rect 460 50 463 54
rect 449 33 453 40
rect 456 -3 460 33
rect 669 13 673 63
rect 685 45 689 50
rect 677 35 681 40
rect 685 -3 689 33
rect 898 11 902 63
rect 912 44 916 50
rect 905 34 909 40
rect 898 6 902 7
rect 918 -3 922 33
rect 1137 0 1153 6
rect -12 -7 1146 -3
rect -13 -64 -9 -60
rect -5 -83 -1 -77
rect 223 -83 227 -77
rect 451 -83 455 -77
rect 678 -83 682 -77
rect 907 -83 911 -77
rect 918 -77 922 -73
rect 1135 -82 1139 -78
rect -18 -102 -13 -98
rect -5 -130 -1 -94
rect 2 -91 6 -87
rect 2 -103 6 -95
rect 210 -102 215 -98
rect 223 -130 227 -94
rect 230 -102 234 -98
rect 438 -102 443 -98
rect 230 -114 234 -106
rect 451 -130 455 -94
rect 458 -103 462 -99
rect 666 -103 671 -99
rect 458 -115 462 -107
rect 678 -130 682 -94
rect 686 -103 690 -99
rect 894 -103 899 -99
rect 686 -115 690 -107
rect 914 -130 918 -94
rect 1122 -103 1127 -99
rect 1135 -130 1139 -94
rect 1142 -130 1146 -7
rect -225 -134 1146 -130
rect 1149 -121 1153 0
rect 686 -167 690 -166
rect 230 -178 234 -177
rect 2 -186 6 -182
rect 230 -186 234 -182
rect 458 -186 462 -173
rect 686 -186 690 -171
rect 918 -179 922 -166
rect -4 -203 4 -199
rect 219 -203 233 -199
rect 447 -203 461 -199
rect 676 -203 688 -199
rect 903 -203 916 -199
rect -4 -232 0 -203
rect 6 -257 10 -213
rect 219 -233 223 -203
rect 228 -224 232 -220
rect 235 -257 238 -213
rect 447 -225 451 -203
rect 456 -223 460 -220
rect 463 -257 466 -213
rect 676 -224 680 -203
rect 684 -222 688 -220
rect 691 -257 694 -213
rect 903 -230 907 -203
rect 912 -221 916 -220
rect 919 -257 922 -213
rect 1149 -247 1153 -127
rect 1157 -21 1161 100
rect 1157 -147 1161 -27
rect 1164 -94 1168 -87
rect 1157 -196 1161 -153
rect 1137 -253 1159 -247
rect -221 -261 1152 -257
rect 1138 -273 1141 -269
rect 221 -298 225 -294
rect 449 -299 453 -296
rect 677 -299 681 -295
rect 905 -299 909 -295
rect 1138 -310 1141 -306
rect 226 -323 234 -319
rect 455 -323 462 -319
rect 221 -376 225 -333
rect 230 -354 234 -323
rect 237 -342 241 -340
rect 448 -376 452 -333
rect 458 -349 462 -323
rect 466 -321 470 -319
rect 680 -323 690 -319
rect 676 -376 680 -333
rect 686 -348 690 -323
rect 693 -320 697 -319
rect 910 -323 916 -319
rect 912 -325 916 -323
rect 920 -320 924 -319
rect 905 -376 909 -333
rect 1133 -357 1137 -323
rect 1148 -329 1152 -261
rect 1144 -333 1152 -329
rect 1148 -376 1152 -333
rect 1155 -367 1159 -253
rect 11 -380 1152 -376
<< m3contact >>
rect -14 62 -10 67
rect 229 50 233 54
rect 221 27 225 31
rect 456 50 460 54
rect 449 29 453 33
rect 685 41 689 45
rect 677 31 681 35
rect 912 40 916 44
rect 905 30 909 34
rect -22 -64 -18 -60
rect 206 -64 210 -60
rect 434 -64 438 -60
rect 662 -64 666 -60
rect 890 -64 894 -60
rect 1118 -64 1122 -60
rect -5 -87 -1 -83
rect 223 -87 227 -83
rect 451 -87 455 -83
rect 678 -87 682 -83
rect 918 -81 922 -77
rect 907 -87 911 -83
rect 1135 -87 1139 -82
rect -22 -102 -18 -98
rect 2 -95 6 -91
rect 206 -102 210 -98
rect 434 -102 438 -98
rect 230 -106 234 -102
rect 662 -103 666 -99
rect 458 -107 462 -103
rect 890 -103 894 -99
rect 686 -107 690 -103
rect 1118 -103 1122 -99
rect 918 -166 922 -162
rect 458 -173 462 -169
rect 2 -182 6 -178
rect 230 -182 234 -178
rect 686 -171 690 -167
rect -4 -236 0 -232
rect 228 -228 232 -224
rect 219 -237 223 -233
rect 447 -229 451 -225
rect 456 -227 460 -223
rect 676 -228 680 -224
rect 684 -226 688 -222
rect 912 -225 916 -221
rect 903 -234 907 -230
rect 1164 -98 1168 -94
rect 1157 -200 1161 -196
rect 1141 -273 1145 -269
rect 221 -294 225 -290
rect 449 -296 453 -292
rect 677 -295 681 -291
rect 905 -295 909 -291
rect 1141 -310 1145 -306
rect 237 -346 241 -342
rect 230 -358 234 -354
rect 466 -325 470 -321
rect 458 -353 462 -349
rect 693 -324 697 -320
rect 920 -324 924 -320
rect 912 -329 916 -325
rect 686 -352 690 -348
<< metal3 >>
rect -14 -10 -10 62
rect 221 20 225 27
rect 229 -10 233 50
rect 449 25 453 29
rect 456 -10 460 50
rect 677 27 681 31
rect 685 -10 689 41
rect 905 26 909 30
rect 912 -10 916 40
rect -14 -14 1159 -10
rect -22 -98 -18 -64
rect -5 -137 -1 -87
rect 2 -99 6 -95
rect 206 -98 210 -64
rect 223 -137 227 -87
rect 434 -98 438 -64
rect 230 -110 234 -106
rect 451 -137 455 -87
rect 662 -99 666 -64
rect 458 -111 462 -107
rect 678 -137 682 -87
rect 890 -99 894 -64
rect 686 -111 690 -107
rect 907 -137 911 -87
rect 918 -86 922 -81
rect 1118 -99 1122 -64
rect 1135 -137 1139 -87
rect 1155 -137 1159 -14
rect 1164 -103 1168 -98
rect -225 -141 1159 -137
rect 2 -178 6 -165
rect 230 -178 234 -162
rect 458 -169 462 -164
rect 686 -167 690 -162
rect 918 -162 922 -158
rect 1157 -205 1161 -200
rect 228 -230 232 -228
rect -4 -260 0 -236
rect 219 -260 223 -237
rect 447 -260 451 -229
rect 456 -229 460 -227
rect 676 -260 680 -228
rect 684 -228 688 -226
rect 912 -228 916 -225
rect 903 -260 907 -234
rect -221 -264 1177 -260
rect 1145 -273 1150 -269
rect 221 -290 225 -284
rect 449 -292 453 -285
rect 677 -291 681 -287
rect 905 -291 909 -284
rect 1145 -310 1164 -306
rect 466 -332 470 -325
rect 693 -333 697 -324
rect 237 -349 241 -346
rect 230 -382 234 -358
rect 458 -382 462 -353
rect 686 -382 690 -352
rect 912 -382 916 -329
rect 920 -335 924 -324
rect 1173 -382 1177 -264
rect -9 -386 1177 -382
<< m4contact >>
rect 221 16 225 20
rect 449 21 453 25
rect 677 23 681 27
rect 905 22 909 26
rect 2 -103 6 -99
rect 230 -114 234 -110
rect 458 -115 462 -111
rect 686 -115 690 -111
rect 918 -90 922 -86
rect 1164 -107 1168 -103
rect 918 -158 922 -154
rect 2 -165 6 -161
rect 230 -162 234 -158
rect 458 -164 462 -160
rect 686 -162 690 -158
rect 1157 -209 1161 -205
rect 228 -234 232 -230
rect 456 -233 460 -229
rect 684 -232 688 -228
rect 912 -232 916 -228
rect 1150 -273 1154 -269
rect 221 -284 225 -280
rect 449 -285 453 -281
rect 677 -287 681 -283
rect 905 -284 909 -280
rect 1164 -310 1168 -306
rect 466 -336 470 -332
rect 693 -337 697 -333
rect 237 -353 241 -349
rect 920 -339 924 -335
<< metal4 >>
rect 2 -161 6 -103
rect 221 -280 225 16
rect 230 -158 234 -114
rect 228 -236 232 -234
rect 449 -281 453 21
rect 458 -160 462 -115
rect 456 -236 460 -233
rect 677 -283 681 23
rect 686 -158 690 -115
rect 684 -234 688 -232
rect 905 -280 909 22
rect 918 -154 922 -90
rect 912 -235 916 -232
rect 1157 -269 1161 -209
rect 1154 -273 1161 -269
rect 1164 -306 1168 -107
rect 237 -392 241 -353
rect 466 -390 470 -336
rect 693 -388 697 -337
rect 920 -390 924 -339
<< m5contact >>
rect 228 -240 232 -236
rect 456 -240 460 -236
rect 684 -238 688 -234
rect 912 -239 916 -235
<< metal5 >>
rect 228 -392 232 -240
rect 456 -390 460 -240
rect 684 -388 688 -238
rect 912 -390 916 -239
use dffsr  dffsr_0
timestamp 1597999042
transform 1 0 38 0 1 3
box -38 -3 184 105
use dffsr  dffsr_1
timestamp 1597999042
transform 1 0 267 0 1 3
box -38 -3 184 105
use dffsr  dffsr_2
timestamp 1597999042
transform 1 0 495 0 1 3
box -38 -3 184 105
use dffsr  dffsr_3
timestamp 1597999042
transform 1 0 723 0 1 3
box -38 -3 184 105
use dffsr  dffsr_4
timestamp 1597999042
transform 1 0 954 0 1 3
box -38 -3 184 105
use dffsr  dffsr_10
timestamp 1597999042
transform -1 0 -40 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_9
timestamp 1597999042
transform -1 0 188 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_8
timestamp 1597999042
transform -1 0 416 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_7
timestamp 1597999042
transform -1 0 644 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_6
timestamp 1597999042
transform -1 0 872 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_5
timestamp 1597999042
transform -1 0 1100 0 1 -124
box -38 -3 184 105
use dffsr  dffsr_11
timestamp 1597999042
transform 1 0 -186 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_12
timestamp 1597999042
transform 1 0 42 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_13
timestamp 1597999042
transform 1 0 270 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_14
timestamp 1597999042
transform 1 0 498 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_15
timestamp 1597999042
transform 1 0 726 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_16
timestamp 1597999042
transform 1 0 954 0 1 -250
box -38 -3 184 105
use dffsr  dffsr_21
timestamp 1597999042
transform -1 0 188 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_20
timestamp 1597999042
transform -1 0 416 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_19
timestamp 1597999042
transform -1 0 644 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_18
timestamp 1597999042
transform -1 0 872 0 1 -370
box -38 -3 184 105
use dffsr  dffsr_17
timestamp 1597999042
transform -1 0 1100 0 1 -370
box -38 -3 184 105
<< labels >>
rlabel metal2 428 -6 428 -6 1 CLK
rlabel metal3 416 -12 416 -12 1 SOC
rlabel metal1 912 103 912 103 5 1
rlabel metal1 909 3 909 3 1 0
rlabel metal1 230 -85 230 -85 1 q9
rlabel metal1 908 54 908 54 1 q4
rlabel metal1 913 -85 913 -85 1 q6
rlabel metal1 684 -86 684 -86 1 q7
rlabel metal1 457 -85 457 -85 1 q8
rlabel metal1 0 -85 0 -85 1 q10
rlabel metal1 -227 -71 -227 -71 3 EOC
rlabel metal1 1148 56 1148 56 1 q5
rlabel metal1 1145 -198 1145 -198 1 D4
rlabel metal1 452 56 452 56 1 q2
rlabel metal1 224 56 224 56 1 q1
rlabel metal1 227 -197 227 -197 1 D0
rlabel metal1 455 -197 455 -197 1 D1
rlabel metal1 683 -197 683 -197 1 D2
rlabel metal1 911 -198 911 -198 1 D3
rlabel metal1 680 56 680 56 1 q3
rlabel metal2 55 -378 55 -378 1 comp
rlabel metal1 2 -317 2 -317 1 D9
rlabel metal1 231 -317 231 -317 1 D8
rlabel metal1 459 -318 459 -318 1 D7
rlabel metal1 687 -317 687 -317 1 D6
rlabel metal1 915 -317 915 -317 1 D5
rlabel metal3 -196 -262 -196 -262 1 SOC
<< end >>
